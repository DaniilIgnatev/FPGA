module top(input logic clk, output logic o1, output logic o2);

assign o1 = clk;
assign o2 = 1;

endmodule
