// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:30 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k6NJ7sKRB7sj/waMZc82ZTqws3Jq3FCjkS8BY/+woY/lR8DwqJ36JR5K8i+un1xo
7N2Xbld6TkYm4IT0lVxN6wAGtPwSy9MgTe/8Ecu3dZEScWXGNxtsiVK+9zPWeKbu
yaufSN/NhjxdhCsWFcp/IV6uFuBp/uljtycrmP4WyWQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22912)
AlyotM6Z7EVMbcD4lDt5rjAG5iieVP8rR9Qg95t4mioMIg3qMkEYhlGS8/VD3pJ4
naM2ysDl3oFrYRqETc8iOlsVwo4KTMaAKen6gpWwJiwG5XV29mgqHZ7nsO3+PoBu
DIq62ga/cSjzO+OtYYx2gOinZdcXmeU1riDj+/V2m5T/5L3Gqu/w4D0b7CQT90GZ
5HkE80/VvqG6ZkEEGJAB/vnNqFf+2uHprmbl43I9XDKDeU6FSjaO+UL9DNFhyokS
sx0RwtJMcHMAAJtLajYeov/4J67o+QK/icVRQs4j2qwGKu2wiKJVXe1+WIJEpWaY
d+wq2S1k6TWpL27NhGELVW3xAf1V1lXlSHBqvP9Xme2LrKA00/h4VUvkfzV34Hly
xnhzVqCoo0Pa6nN04Bgs3/3Vv+Awo2BldGnkDdX1HuIMY2SK9rtrpXKM7fDV0Dmx
UFhzN0EFuydbn2E99eDZkFY4N0w/kMBqMvWqZt9Iii7ACWBMom8Ijj1B/REJX2o1
RhIaYXvOklG7sUvBCXC1J9viEL1hqibWZTm72YuahLiLEa6cDKegiEVih93KusrV
+jHETgIxT8Rh/x7frtFY8P+5x+X8sJWkib8V3WF8BeNFebRmwwJK5Br8PyQVKJqG
6aU/5UwzBhoGUhHm7niDxnG5L15VHl0PAdmVfQ5rVZ3Iac8EBpnUyfN7/RU/B3Ev
0RJaWD+pHV5HqVng0dAphMekOyCzCIins6Lpd2wnhPswRxyoXvKI9ZbubKB8IIcb
Pt6WBIjcvBShN3tFnS0O4Rcj46oXM41LfdeT4Bul00npE06AL7WWplkYGNBL1cjt
1XmJmsi6qO7YrmCo/272tYXIV2peKZozvGUADmqM5qTVU+GCZqsZyfbmYieyXS/N
8bOjoj83ydzwBlCVtcnQ9OUk4jNnO17C0Pgn/sURKmfYVAYBMAAC2l5+xofh68hM
AGtuul8lol5GNlZxPLmJt0aGiLjwH9/NsklJHtgnhXQIv2St2L/XPIHf/zePztLo
HegYEnERPx8T9Ss/2SBpw4FP1pziNg6DWHd+nyXQtEG8Pfx82m6LkN1HpZ6Nt21x
qZ2AyOi+Z5HhzamAh6fFBvYlfDXyINU7zV2QSrS/BkvV+RDwpL3Fku6od8Jog85+
vPlKFdOyBJ68aczaKnOePPCA8paVhWF5ucMbAxucgXuzYTgjpvfFXX0RZ1d8M8Lo
N/RFvVbwxs4tAd/c9JtUlVnBIbSEAnLSUSA/y+SEIJHNJqvYp7HYNI5nT7fpOVwv
cXKwdvV4RBLciD2sNB1lyeExX2S7tbEhy/UiSwVVmHtZRtieZ1l7EvCiO49HYNOX
Dk5fnw48Ty2n2DHqnPdKvFDEiWtvuOXksE41V30ulqDDkxf4M5WsqOvvaF1ZVV+s
jy5Wp8zPBYhNUkWo+ZK4ekjqgy+oiDHkwo+rRN0pgpMENtASEuiIagFWg31XbtPd
LvWI+D+XAKztulWfPP6SKcNEwswZHZTQfDI28N69Rv3tIK9ypphABpy7zJBx2dyZ
1mBZzWTu1pr9/vgaTuT7SyZC0Ebe1iwbjb/2DEbTET0GMVyg9vSMPQxZmvGTul7/
DBPs+u0Fip5cSKPxkbGyWZSNlnA/bkPC7bJzpzkW7CEB3BJ9nvc36xeGD914t1/r
J6P0LFM/VTa19tWmBORJB9AFsyza1zygAu4816rYaQ/TE58uBBCKoczvSWjOZcPe
nVfdjIsj6zKKRWh0Ipmb5YzazbwhZT0bpdrmW76xokB/4yF5q2bLaYuDRTXyyJYe
Gu7FUvdAP5W0VtjXcziumxOooMC7mZkyFeGHDt1NCsF/dDR+AR4X64b8CYfiKWQi
NPcdzlT6LtwETyGQ4W8NgTrab/QN5PX0xjsnS7e/GuYOpExGFTwloc7DCBTWNrjH
J678QE8s/gDa3qJE30AaqY4laH73mS3LEV6bRDRf705ceuBfWDxZ1ls4wL8SdvoM
CLjpBYhfw4xTUI1SjotJtJLK1oOsYRF9LLjMCOQBUvzgOQG39Zu9gIS5UMx/QbMG
MzICVGcbj7/mikCSUbz21aA2DoDBPyUYmqt+Umkx9/cfJ3NQbtAQQ+4k5VOpAKai
kT48ZQ8nEVOk7xAhvYFofrBqd7DXVYCo6dClEJtqqSKGCcBDqkcyGYd/yBcOY8w+
bCXPj2GGNkE5H59ntfY6udNekM/hWk96uk09P7J57L3S7ho5h5uVZDbXxNKEJLaO
wAU2ChFyNflDDk2X2Z9ItIMHk6qh4x4r+c47jdipK66smx21Cqevn9Fqzs9dtOwO
r5DV1Dhfxi/tNFwBT977oBuX6L555rMjv++J+ZHySiQzgOf2C7z2ZHAJK/h4WJ5s
NtN4kQFMqfyhPk9J/djQZ5uPJyfXJVnGYsoVFdlYvyIvOu8ofhWgszE0CjD5GAVU
DWc0S/gq8j3oAENjBQjoPruGYeKc9jdJ97dNFHkTHcINYjfQQuxQg3FSfHminJPP
D6BxmMui1vIeX16z04mezQsUctcuH1RQHKP5zxwG1h4js8c62QAXODdTAZnm7T5M
gMJ8+KeYHJhUaMB878ZavIz7UAfkiFPry+XvStApEDGP3ZjVds+FHnvNT2LqKENm
BRclxLmvqOymu9NoAa/XA9wMdjK/Rh+z3YIRD327+5Kc5dunye7xxdA+IyqtiRdm
/f4DARphNFI46imB/uQJLczFS8ubB8ueh4gnAjB7FiUSclcqIevQYIc/H/JrVY6e
X2EdTf4BlCDrb1JZ/FX+Tl7z1NuEiWbtHw2Pwae36mdAHQMBIdV1KVnTaxJx//lq
GaAY4DacDWNiBm3TnK9hhDXjzHMSpvz3oT8HMZaKI++APLFe68AfGpApuIq9E+bt
/Xr4JjcGVoJF93ZqiTQn7OJHWEjsdaTeLD6CwHirR9+8BtEocgR6zsxOiT1qkCVN
23KyKuAOxsQD0TIlTJhe7l6VnSinDpWiMq6h/FSgwDxiNoIcDBMcgIksACjaqqJK
LCCRwMkSz1hS2iexmXFUX/deT39vI4CzNgGLzKw3w6Rnl2C57g5SjmtQgcH3JViG
OoSRnwgsmurAlloI193GeLFGB8ZgZNZp87EmDfqED6rgizoQxWZ8QZ5bqEvXOOOD
bx/sNWF8cCsmk5qkhTwfyCaAyw7xo2vO5gysC/idrO7QqsOK3uc5RoAnQtN5fRaf
AvCU5+XnWwuIDBvgZE9WPdfPIDxIEcah5m/sGe7jbqu5fmxqPTeOIn6uZkuCohzy
WNaLRh5oWMswoWxvFoDflrBAPTdgeQmaioKO7VPto4wTPynyovDhqoj6GpldImlo
9ahKh76IvCo+eL7zHhym6W9WzmhMLM9flNwSiI5jr0UpjDTFruhfS7Fcn9ejemvN
MwalglDQwzTVeZ3EqoHyccnbLd3KZpQ4HrYOasDIKZysv2laSKtJoJ+nN47pRQBO
xx1El9/d1gQ3xSTXfXtkMN8m4TRcMIeYVaeJH7fOs0+/wJ/guy6cpxx3w9rzbMhi
Anu2cQhhaxkiegR40+zNwftHDVDrIVQiqRSGN9XBz88BpH1UuKHidFrb8Abwb+J0
/qEwqq1UV0fHmg1EejfxvDdxphaezRxGAGye+3hmUzTiAvqfSNBMZEgBiiVE14Gy
0c9eLgtSLA8ccyg4d2SxEZjgFSGX2ocF2/5QHSDlwRtdOa0i/bM/eKhzLD0HstlF
J87X+YYDyXTRF5dLe+GEnZ361DbkmuW/OjbNJKiiqVKZdWdBiI3GGiuOEf6ewNaI
K880nLhOiVJwUb76ChGHz0wEpDwPnP3GwJmxtuQ0/zuHL1RNSq/TKpip/1Csu7Q4
JZd9GmR08MWArGvICQ/kNFLZDcsBteh3wDnpA3J1oQ6pdmG8+i8awO0mzOvnPHhd
Vl/3UCgsV/nFl3KckFsYmuCW+L+fcZ9qdRLzpKVhe20OFd8OsVtUnWFF8LyxOPZd
1ymIbnSGjQN9gCKbY09m5+pLRDqa6a5Jcql2lqDqlcjUcPzhB4SqTMK3hfZJhMv6
4vocN09lYVrLzd5G9WZiK8xKEd073lnQr1Flfx0Ury6FiOmphzEl+s7jG0GyWHDk
1EQoOlwFM9MlDNspOXYk222OIuTYo5/R747adyS4RP61dbFg+fbz9DCBiS6kPceU
2pElOU6aAzrGvxCtRvuELzaeGOzPPikAeD1ScX4MvfNRx914hzkxa9vsoKBntyhi
JRu5EyS1Clq45/zuWMlyZkVIiRsWQiPI2EV4M/5ojV3KvoEogsJaGou+TlFR4M6G
8mwTBAJ4S1Arv42gqNjOibn8TD2evJk6XBl9Xsl/PglpX/ubkxjFVY38YIhoL8Z6
XXgNCWPaSOH8EmulAfsFKI/pzDTXbS1wbAI2tn6M0QZH2qiWcLPYBxE9e3iifF88
sR864Lxgv6DlIVJwg7FnnFyTndMyQoUTLVgm690vcyfDZBzpoT8XXarQH5v5D2ra
w5x4xtnbRTjfQ8Zzjl9PvrO+0W7h7pNKi72DplJlOwru+Zgvh93ELmooO+VLMj96
C+6WPChE1vegaF+JNJKcLOrBUx8Toso+3xEdARGWY/YlobMJCfY31uo/GebRjrwg
IyzVmR06VfUBCnSwrI0iZH2VOywieyspP2DBfBhO5plV2HQ0pTzW2CMaIPwBUlzM
ffDT+wkPpoMUrQStmuK9Q1xnSk03KV/vIwuG7WkvjTbpTowXhGHTOLRL2jlXtMz1
WmqrTqG7iIG2cZUiqSWu6tUhFZC+Vy2NrTr54Pi8q3HA1OrQ+dO6U//gQXfRq1vd
eG7qvgIZG4oRt4oKC4Mb0rAUh2cEWFshPIPScItO7cSvZM0Zm64i2Alhu/Gfmxle
VU7YY7Wjx8T9Ieufe47eF0JGazD55Yfoxm+Jwdy7pgkHvebU4WHz9lqcnntAIycL
XovgxTFQlVVAAorQSi+2R3/nhyunrtBaXBpUiTzWKcxpOwYbiCHplLH2J9HefbZZ
Y7l/ZqUo8/eOwGoUohP3aP2PTfHY7/FF/LLloi9KdaalJCqsEaV8X6yFr7SuqURX
Wik7uKHNnzi+FngZh/EjN6XjXEvzG8a8QZ4A1nkdhDfoeZRJ+BvdCryhlRaMgnS2
bd+qZ/O1FT4pNB1v8z2z+73ah6Wgwb0YGQ+xAvvpTAT9rdDG6n1F6y2xoao4yKTA
/TzJasPATy/q8J5Xi5BtvoCiswwbPL7iUQL56i1O0W9JZMI9oQRCa5poM/aDuQ1i
tsWQv9I7hCcYpnAyICg7NsLS8lPqpXRQ/l6Cq9C3IdYkBLVgM7+nXm37mt6VCosg
VQQMgKQB1N+0mDJMHvrNQXdRnNu1MD7eBKAKWd2z5bA00yrdl3h6XRAgjC26ndFo
xIdDH5v75vVbimMmNz9Ifw2xsPWsTAW6W/HUskhmb9UzbnJKZ5hlHW8LWK729Lwa
V9DnnSzwVQ3/WflLK/wBbi8nEsEA+lX+JNCxR2lVoSXKRnPzSDPMaPP3eTr59TZI
CTfo9Odh6vvHrfSWRWgmyyF4nS+Hd1Nev0lCBpXvI7AikUMOeRGmOyo8oUBIG5YM
ZIwEXM3a4daRUluFJM25TKU4MqCJY4KqoyTWlSvvjDGAtO8IUp0dRChRocU46wGh
tRws/UaE57iCWB9F+WhJQC7QoutyERkwKJ81tayJrMbcaWnIOTbQvj/VG/Jd4EqC
ZYb1rN6hFnetbgGbADOKPLnFVjEa0/mgEhb+6/brjXVXZlYulr867h3z2Rcd1NCF
OyQG5yMkbVSVGNPCYgbboELaXCXgjS8Y2laZwPip8hWqz6nf5/x+/Z+FkxwNNwG4
AChqi1r3hm1MlvIkFgAJYm0sp2xaLxSehLpdKCFcte8u1ccx6vCV1Q6D7TSd5LuV
jLgry4HWiAro6AE3nQ/rXtro24RmnPZiX19Lq0hgr65b+MUOc8lR2mYHrri6Xbko
HAfTroF2J4MqDzb4gQX1i7C09gsxjbPjtdVVhDXY5+nAWw7ruz65zM9z5I9haYTe
ef+PJzBEIEvOBlfj1t9gdqQCz1VhqXaajD7IdsqH85Bt1OP5jBrpKhxPnMLCBEEl
nZfCJIJH2GkL/UGPEeUzyHfi5SwZkGxQK1IMvp0S07J1ch7ws8XlIwVcJXkT6AKd
S4yrjQXLPh/0DrIeGHDx+OJADu10qu01rdcHHpGdSyMY2s7/Ffrxn4epD2dEl1ZL
T3NdNavOEd0/YnSHT4VELAlbZJG4zV4nAFIlpVHkeLqawTlOYmCi0VojsC8R2umP
eCTZ0c5YbmHUMXAOTj7b+jzTf/9D6xiURBp2rxpLG80bnrPqTxH3BbCgvvUWmMLS
Sq/jHGOmsAY3yMAC/FGrC2FWhi90Ov5+C1/UwXIPtLJX9/ZSsQE5pyYtihPy+8q1
3/AX4iAIme4jIl1FeC9CBOSwT87Rv1Ov/5YwRjwIpC1usnqjO49e+LWxTt0ZBGQg
1tNJ5a1gdtDXPf9YSjAwUmhoOdP/4NkuKcmPZPuzPx+nd3BYrozQ7GyO7kigNgh8
1PL/ihU86I2NeVFZJd31Z3YIfMc3sYd3oaUs29oOtvXnY2xgCD9vYvQDnsmt2RQX
mCmwkaD4oLSNcDZRzdM3Ymjtwn5aTa7yPrQIzQhYDm+tGnsB+rlj/5hohi7oS07b
p2RoYLD4zLGjHr4S+622BffEGnv+yw4z3qhqC9wxA2PQF/E/Qjoy8cfBkoAWHt4h
IBNU+m0wJw7EZXP1z4NFuijWlHVaxfw5wSGv3vN6b5xsXgAY4W11S+LB6kiXWXju
Om4JvXDKJfgbhAgK50Crv0MWS9zNGCw2yVkpOpZ9IY4NEPP/oJ08yBXjw4uf7tzL
jPqH8kDjKIkg/jIZM2uJYoCkjtCLO4ni2q00ZJXEKJGhitux2zOmSrclxM2rXs5v
RYVSK83I07Dd9TMHx4FEwvDOugmR0kxAuLx8NSRA9t+JCmBunhrPsQBL+WosCAys
zXCNuU4aJZ3HPCIZuTXSWXlmJJLe1KGK4JIqfKJtMKJFBalRg7z2qoq2xhDR6asK
dlplvvc37sZdI7tgBSuoPtWDNhb4zMltjfxVbrEoP0FXIUs2lcREK67YA5S0o/Qm
+JxJrc2jqFiZlGKc6Yms8Smw3tQrxI05i4QWz7zOfPM/QAB6dd8EmPREtXqu4PXx
Hxt9nyBJr558bX4b6x12exqed4pMbOZ1mKguaxhp6NaUhZDFKgQpmG+AZyeO39DX
A6jVBpULW81wE32Y1OdVsSLWutx7VTBzgv8+q7HYvAw/1ScVn5Lzj/dw8WURA7aI
z+qAJGNb//eB0zT5TGI94to2a4Dlp4/L27SgInmbn7+UUUYUKI+Jm53DTqzgBGRW
FYP8r53FATzYBX5jOSNISRSM9DWRIAQMTgR/78yR3AuKJuDFTeBXa1wnuh7bderv
T1Xx7zcInryod26wg3yUITCQ3gq5f8nPhG7PHk1ENJ//LwLUbZz2C65kGEtPJY85
ScKxQjiIT4/fp25zwJo/fh57slC6b8YxikrQEMf8IaXKguxD+FyXVChMo20YZklw
HtrmjfB/aoLCUE68Ot+fm0+T4CCaklIZVRUVNK0UtL94yo2WJuJWTki5aLlXO7aX
HKMBAfWmJY1+/JbZJbc8rRsb4qZVOHopWRMR0oP9VzEC8p0uYUHiWxqlwO4Zj1YL
fU0YOEjQ54Tz6WmCaPnGEC/Ut725EUsK5Fh5YlnxZdvgYvTUwpg0g21rmdpnO32u
sCbvrcpA8gJPuVtIMKIP/NVkenuwJduTd+RHZpB27LNvK9iwG+zWvm9FrPmOhvvZ
+6NIkwVY+uPb/ulnL8POcTgw8mc3xeVxIGw0Uum1z+M8p95fNOOW9Vs+aNsWonXf
p3WSEVZwDMm257WOQF8jY09i6mxlPL4Fw9RlAtpDdkTjn25Lgf4PkALfxZkXxfzT
7YOit00nYbrCQJr02azmXGAolHtslh6Vu2kCCBYOepCC+2JGp6wQoUEYs4YMOSGk
d0+KHpRJmNcSV/zF+lBiGiElV6w9uXzWDa+J3K/P/09J8zsrZycKdK0aVvyTCBDs
JJCpSYRxbXKgz5tq5Yc3W4wAxQV1S+jIPESkTDZRCKDhf3d/GdIDBa5Aqy7RjwtD
ILVKm2yaX5VrA6TiKdH1Alzmpnu2bvNLMTmlzOIycYKQLk00UVEpoG8ut60CqITb
l3pHdOQY00rzzqeMjWQ/HqVCaKLffooRaAOyu163B37PX61dAtdu+Nv2W8Ad65Zc
5RFG3OdTIhvG4NMj9+POvqduaWLmVA7as2eN2quV3Y7ho1/gPWl1zR8A4vMSeeMe
6V8p+/P36jefNLzm74dTzxA4UQLUUYbzqnIhK6XkO+78mCENBQUYMt3KFHEWKir/
hFJPjgh7xwnEtLkcACRKKji8kg3k2xYMJrbEWi/a2ffepB6Y0GnqFBoWOr5e7AQO
C56wMhiScLIUtRqNC28dnTRM8WdKkoPWHcQTMCkjsuGGan04KJwNA4MsZYy6oyhE
6FebaP2joX7cJkRHYpssOiC0zKXkEpv+FeIQOlitC8QSKuQAvx1+OWqt8PVM18NF
hmIFct4wpgeE/M20P53gkm5gInZLg8u87DFe99xfRvePV8gPVJQjm4Qa0ylHyzvE
BnG3sG6adgS7snPmfBg1eIGVlwqQfam80I51MiFgjhqKBOqm02fdx/8qcJEri+0v
SUv7v3X0L+IPjyCbVRkNZVKKzPSNRSRHj+MmWcmX0VSfjiqB9N/zXIIAglXE6Rz1
kxtToO6TGJ4UCYlOzc17l7zVsWz1Fr5iTY4Bt7ALyxCW7ciztcSLjthAipqqENuG
deM0B6Ijvs0y4bwqPgK3dabquRBTrvEJT98eacdo0Eooy/w1Jmae/U8LtNBkt1aR
g3KWzV7zGWGbHzaETJ4upF/KQOaoh7W03OGkTsApvrGXbUdmB3VbClwXFOzvOzjU
HcwQZfRdvrTZEoJgW0eFXFcpBn9CUVCu7mIpkvwDGzfyl58qOa04hK2bpmx8+mNS
dSbsNNBTfAUU81ITJfNoRaBhxc9BgxGOhBLk24LKQ+DhzTcOeiIcS7zrKYwHBqq4
xoEOC9NjY4+5KkX3d7Z9VR8ML5YugEQQT1IPE4zQBDLDolwyiRSQDy2U2yqsaoRj
E+4I2YKZAyoWtLo7DZP+J/Y9V0Cj2WuDaJGEoeTxKSDIZ/ijnDykFjyD2YFdjD/V
wi+mFOKrHfbtwMBQ1kslK6ZPhqB7BlXah+yRgsXnRJ/iQYDQwZvI1md51F1GCWXL
rDLEV4v64Jpltwre5gMacPDIdSJ3OV7pODtc70J6c8GMwFvC7hNzeiI1Oiyu3t04
e3CeiFvDqaut08WyqTbKDDTF8l/IVI1hDm4NEhcce2qukP8Ntl6knj/FL7SNk99T
A5DjUY77htZ3WWWjvd4iOp/kXUAE/B1QQfuOkuXVGiPD1TLeXb2HmmKNoIE8/BSX
YI+AJIc1vyojyt9LMWxIy7Fd8FrQRuTIOA8nHuEnRThc8D7acRmtRni3la10hg9X
GPa7XWlEYsGsvVAvsC0NnuHm8xiLTZWsJtWLx3L8e3TOqU6tD7MsFEzVP3/sobg2
gaf2YHz7AtwgBaCSuAfYVZcD4GgHEyhCPjngIGAdLANmgA5akhvx0pRnNMlBHVwe
QIhdxYqkl9eNw0qsbBS+IshxIOlHfcDMrVA+zN03VA5FoFpQwc3EcyxVEvo0tTSQ
iosvfhZC1wAyCc92fCT4nZntt87tKsaDqq/umXEofrBjZQwRWFXQIhKTG4ZYrD2N
NTQaezeaTPrPLZxuNGXWyPdu5cNomLTABojD1e5k5/Es9LihxxIpwV6M5g2yfC6P
c0IweEbJcdz5+5djKY8vhltLt4IM9jBbtKZSC/2iBS6cl+W8c66yakTdOybFw/ej
blu0eahBR0kYj3RxY92qEb8t8QDkEOeT4hHqJHYkUtOUm4Cd9cnQJU6yYvpIKShE
Z4b1E/hz0h+YCikrAwfLw1wKe2PIRC67w2zrN6LxEYIzto6wurejjxbf9DBFZY1q
xrQjv92ne23UmcCgHxui8+Nco13TC0jFTYEEcKXXTDdkRhggCnrZwH9uEgJhCtcc
yQQ/I7nN4GCq+vwhBcWihCaTudU6arm9IckHkx2KOBlq2aMbCAZm6VDwRPxcFjQ1
k7qgtDXkqyl6NHhAom7oyc41NFAcpxbEoPk5o5yhNCJCT7G/7ctyZ+c/xqGBdScH
3gLJSt/HwDhdGAFDVXiedR1a1IQu92v3VZmoZBkfKretu5z8aoj0MdhOuAGV2y6F
CJ+WM6V+lHXHfL2Ab/dqbTI2rA7m65PhCpQLzPT+ZGcPhftIey1UGlvLtXP7wNAQ
ulO1Rw5Of4d5LPsnSaOZdeM1BfnFtAIqzJ+ihP5ADS1QwWcc6W0nhcb5wk1q4DQ6
wBJpFd7XRrFU6NKlIvxka5TSf5H5Gw3C0/B5H9ZfCchJcUormvwQw4rKR+zT5aYC
2Ao5wTsrPLpVA0ZAjnm/5JIUaiXBHB9B6xiaoooKHvKfeg5/TPhYaGB8Yl9UB5zB
fkWMPlhunzWfg+RfhAHZIA9SRhgWEXAliLbdbQ67vFS6UwofFU4JoAg8rZ0lqh9k
lxttXYuWQ4f3bXMyDzQhJPdhmMlpRm8YKGrw1fVnfLMDtAQIHt6XpdXD7kM+rNE4
IwUZ6/hr4ZAkXBlT0COp1LBGdHA+c1z8cDWKyN4PyffZTYNYGJWWVBRMOAaZBr8d
zHuQsLNeFLiPPjk75ikhoemlWhxWD6I9zJ/MQ5Ec1hjN8gOK7eNyiTmbRsTA31Bt
xsQ72bGP3OOcWYdQ6h0Cfeh9Ypmn1dBBaQxzXNt2qvFH6rtv2rN7ki30Sm9egr2Y
7wYEZAbYHR0naombp8nAXSBHr/DisQpi7m7aXw9OAJknecsMiITmOP/G5oKI9gTM
EuXt1+RvXcSrHSc4155Y8Phjpef/Bc7HvAYAPX7MYiFv9y+AZil1lb3Hmx6/pbUT
NPHYx1+oUGvYgZZMf8jjnRcF2a88uQzlecjv0f/iiixUQ9dZRqYfyLM3cQB9ibZ3
Gku6esSi5v49nzCTf1kpRHFQgqmqpPXi/X9Nkj86c70cM7m5baNEHyQ/x/0SytJB
dUD7tTUpcXl0QTjt/Jp/FZ7lri2Hu9VGVECugFCp+jviiF4XmeePaRZ0FTRdG0qk
7rGcWdEZV2Rk5OHlJtnnbfYDza08ZxU0w5Q1aIlWkweSd8/3cmbEC8g6ZkfFqQct
Mck8EGCvE0L+2zdTL+hFTTTBXxVb1DUecMFbvVgbOz2uQs6hPuXRQ5V9xYY0IdQH
BXNiqjbpYbfEM0TJ+6mtjm5/OKXHVheqO4IHMweOPMHTN1PfColmCilpMjeEElEP
00TkjrXLrCoU8FQH4/NYaoJD+DhEzl5m1Ejr46Jn+MFnhmj4t/O0E2/2lBXAIdfe
fzBzy8WmLWRaEfk37rahsddv67onD2b4hNdFpKqJNlTlN2VcSsTqPasPCm18yHB3
2bcdhxeGMr//QhM9zzTHCZ0aJQbIzdeM1VFxrYH8vpYDebyx2QnrTc03ZDHYvPfz
8PG7vC5fN/+8axe2i3u0O8nW5tTl6w9NWaWDC6a+Sev+eLGZc1fV6Jo6gRJ1vkpM
Tgmt2OIe/OgYnkiBAmu54et6q9pgR2MoFtH2ljM7V1+Gqqe+Jjn96/E+8j1XqUTW
h7jnaCzq5r5aIDkNvogoIL3tn6bH6GuYnn2O2EoKFVgyzDPIgLSjkgtt6oo8Cz5d
7ig9xynhFxkJmOrZfBYncmD8eq+W92PfM0iV+HP15NJLPvglToUQLM9Iu47MZrRU
XRHdvLREvyoRT5xDv+c67slJnb6t3Afs99wJ6v5xuuBzCNMHKeWFKoYKQjGvkVbP
ybz43fpFiCaoD6LMO52o8cMvp9CyPndNa0uGeX1IeZGoFF3lX5Uv5OQB/UsAkIvk
oPrrYRZR3Ei6RBj3On/PrsMS8h/qoWXSHRmGSI1crdjuQM+wCe+XQU1iizOn/iTr
Riip9iX2lvom8Mrp/PYgnFk5uaZOl12aMO0zZw7/tTp66nz5EbC3VWQEqEyfNUIp
BjVdb5J44EcDu1K/+z3CNvMdpGAlyOq6pD2cW+I3rrRNg8a4aAaLgL3kb2CGcQIK
IsRjzRh+WGY7nsKJKYNcUCCq1wmwsmNedkexoVZeXSoos2gr5exkol02P94gI+gn
lnuQd4BSNdlcP9VZWlMIfnHmGeenRtGQ3KtICWSuVOr8SCZ9orXUoiNIQz0sglc1
r0K7w0tgXUBZdcDTGjv8b6DNv/xCmxp1Dwa36o47ZHnUNvjrOYE2T110Om8AnvKn
gZ8YMcXnao8yGa04P2RzYlLDXjTi685S9q/4dwpVYrk2jWzu2jUKyREfhewBFHP/
xb79WGBWoAvH1i/Mfxgn7Fccmk3DE38pufGRHpbRtAlPokQS2l7+MgCFI3LhjHm5
xZbmGBHm+GitQWwMyNjS2ZT/FsGD1hIaPSoTCv6/NoAYsK7pWTYLvcPT0aQbRSHq
1U2jNJtX9rhIHNPWB2lEZRhvq9TR97xKXq2++48k2palebNMzE+VUljPeICc4KFp
u3BujJuuHygMt2l9atdD5jUsPlfKb8uqwKx86zaKumfgMhGsyfDSyUNR5pw+iSQ5
uCrYFrm5RWC9vMKL0x/0foCGDFfnsj/nPVFoyInxzKwxhx6WbyxQYvlxbqE2QXhE
KvxzO3OEW9ppjsJ7coCj1QrTTWhz9AIQsCRdOnORP+Qznps7Hv8widcU0oj9nZLm
5hLDUyXY7lZjYcjZF6CKtRmy0OZjbxJ/feXsCQpT4mMkGeLLHoLRHXzzHLYuFgMn
qPpbB4/LOjS1Ai+6dfHEa9fw1lVmLiTgAnG8ZJ+AwCGVYijLUEGfkG8/+Ol54b1b
1MyVW5gV8JUXYvrJdzLzEIYM3i7pmzsbdWmMUgDmpP+T8IcGW35zBMTvLRdecoDl
c7AM8n+q815s7iNB8RVd4S1UWa8CE16uQGyUKMI2pY6YKgz/lV738DjbvGV3GfFQ
m+8d1vqaRGsSPylyIF7IKkyZOotEnGytQL+0i/gc6FccikUwm2cNbh6csJa/8xRF
hBG+lCuVDD359NoIr+5New35LDL+TqfF+081hvb76CVhmQjjxWebm5XOhIRVHIok
Ya5FhGOPuTNp3y3qqPSjoZYcILa1jvKB1n8zsqTmk8ciC9TZBrKk8PPOsx+F/1Bm
u5kNh7tEtWUlml1kSM4P1B3BXQvp15lp4ZylFPpb2lbIdgpjsYY2bWrCEAGbT56v
SRZL5CXdq5N5H9aNZXXD08x4TgSUf3Bm/+76nhrIJfBUlup6/ZCg2fGksGoHfDhH
Et/522kA7yjsE8AaXcUFwdFUpVfbgSf3lNnGL4YN0S3NteBQUNI2wS2ic/nMeuif
xWHR5kRwmTJ7EtR47UNpol5BnH6p7WyuKQar2USAb0Rd3+YQVG9mUHOGQgOBFOx7
w723QPeU6uDnrGoaia0tG4hn2QkojpfqstIPMICahS4QRSkDduaxEjWk2/Zfbp7e
rilJEZl6hEVXoku3zjocWdmnojyilo7B8qn/LVag0jT4zd5BcGpgzAzM7qeVsArK
DaVb5rlbhmqDwHCqaTo6hRpmHk5UeCt1+ML1NvhNVrh1qqx/T/OJMCpWda1GxV4D
DafyRGzGFYHLfjkiC1BDZcEl/100GCWrGsCItphuof2jn/pC9HV7JUO/9D9THv1v
MJl0NMJ7acxEbTtqGHCiEK7AKVXJv4XndVTHV5dJQd8ThMW8iX5qfrHbZKg7ge5S
MF8uMM764VOcDDX9+BPDNYfBqxvgGLzG50+EK5aqHS8aAiiHJ+WfgqpuQJFP4YEe
KdvXiyft1dtUL4XliJujVGi/zE+cDerD+nwrMedgw7eaCR09Wz50nVaxLKFloOdb
Epsar2y9s1/TYQMon2KV2NRVKC1AJYXOSLGkghQjMt7XBuhVqekLcKz2CJ8sOE8V
3GZGRPesEQn16p9mNUi/Yznrem6xP96CaTltyuy9d8pdM9pvtYuE7UatfEBxn21Q
m9VzLmidvB8WKrdfMmqyqh0UqCMOTKXuLli37QGKutKCy6veduqeI0HdsqmmyDue
4rQeZ0cQ0ZGYSmRwsYFTBDuKLKPQ3SAJ5FJr1os3FkyqBVXtCgw5ODdw+eYklqX1
COZbT3DxhkykPkrMboZhvK6I7+paKvZVl+XaHRlwg0t7KLkd+GbHqfNix0Hku2e9
SKE4iGoEJeSrZx22VOnsPfXr2YcBuD4+bzn3+IMamDgrsnkYzJyqeP9/JlfuieY+
QuzQKoVYbKPmeSIpTRW5+RytRJ/ziqtVKjwOexbY+p8NRZEB3ChPSRp+2ocipH/m
5tptVEBJUajWucz/T/g/wXqA6S6diFElkwLxmtZVELcpWlW9NgFIOIiyYN/VD6eb
AyPNHXmO/wJokxbAJ7FyX0a1dc9oMb8KnAaKYlkzkbPsgNA2bkwq0qrax6YFcjBI
3kbgnb+fPVAgdDblnt2cgMhl7Zp9VNzlw/pnS4/tlhgCMIvUcYgI/n+RsuXndMOG
jNtui/1RZjL3SjmtPd9c2SaNUUES/saJImGIVE3LU3UVaT0+95urdH1slkZCvnTg
rKHoJkl66r3h8t1Rz9Z2sX4rKkXb1EzeGC//+IAArDVpDX3TuU2uC5Go/j9MAofz
MN+9oUZrrrOUOD3xJjVliAoweLtCTilLNXF/Gl+kC7PpfGV3MTnOkzVmfOkRm9zc
tvdBz9ntHwyy1Z3zdslNyICKCkZ4ZVr3XI6xhAhIoLrdCbthrVaUSH224yjDwPTl
uIpxOrVgma6pU5ToJZatDiLjQeufMO+xo2QhQZ21Rt+KMr0PTFtzhUnxPOnx2fiK
xox3A44HucmvTFznp5z5fPxI2IoDUTzWhKr704TdaxZ/B9hz7bOWbT7FLRIV/Sjy
NTghhgzolV9ekJe52Ka+bQnq/i+HY8JXBb0WhDGz3YaKQ9Log1jpic/Jm6vTUIpm
WzaisaKQ0NndSRy5qln7eCKZRqh61RfWWBQEKp6Z774XqzTuYaTdSDSxCwWG8SyU
coJ27Ejpv6K93ri438nc8MLaq3lSx/+mWHdOaPlm0m51XsfloAbveOSd0yxVYgkt
4Dq/l+Cv/Ik+FAD7K/k4kJWst7zmMRlWXKIQvMUwsN2+LxsZBXuz2oxpmqlWfDZS
qSC+L/3fX8D4k8GVR87dUKU4O81AXATrPwfzc4REOXu2FlYrYGDdePiHwk8GA0H5
uqbxvQldDX1/Wqa4UvcsIhIUvg+pJ37oiPI0CyzJz6wY2YLbgjKHXrduwK/3QZme
MBzxAaOVbfH4rVuYvaD6sinDCwSFqXtSdy4TxFs60v6QWO6trUGGJ5J1f2AwGtsf
y8dXwBD1fNck9Yc4wQclZdIIoqjl71pEhxekNHcZrPXnP5zjbWGjzUWyCHDWREYG
LNi5PQacyqg54wO41UeqJl3QnJyiRD7nk8K9IgO6lpbbgiYpPkYe6NsOI7tHph5a
tkCYSK0NQw+mU77s1bLsjY/UJg2AcZEqfNoGUL6RDCdB2rqywoCpQOlfwMmg9RfJ
jn7eGnE8tDrfVwGSfVSIxxidcpe57NLBe9uewN03O3yNTr3wK2IYf9V/BjbFu+4O
x4xFmDVyuV+BL8MX77tsuQL3Dh9Z5y1fe/Srv3ST7/1nYfHoyRhkPwnbaVyqiS5L
oWLp0GM80IQkwsR6VgQPcSFeeJWDKRi8ZSRTKeeklFe7YhQZkgSF3AbmaadZmzCU
YtCjJqKIW2OejuWKWpgbQt2+cFtemiO3l2Wbae4VovJ9cEL6Wm6rN4rAZQl5p1mS
faqyp1ZUqPWc2V5FOi8i5EfNAlA1PWO5eO+pfHazWA+4jCZpmZXVzaiFvIH4oqoV
Zk8ar9rDQNkrkbaTwwMYvXE1O0wR2edat9a9dIprAOF5dK81QUDJaJ127Z5f9pa9
veDO5U98tMU28C3Qmsdck9lAcpot9FJlaueozEwE4rfTIxcNOkpb+cmR9AOftNMr
0cfZrpzfKCt3Guj2gxiQbZZTsKzwH9rPUaC1RQi6064lBWh/LNjRHLLsn7grimru
g2JAWKR6KhQe536g/mmN/jDcAH9alA3EUxiSyWKTVo2reX1EMd2UY34OeMC0hKy/
iSuYIXAwzUXg9sHHNI6+HFykt+3Ygykj9w//KUctdfIxADerLYFBKKYoiM3TVBFC
NMwIDZCZxx+6LBbMhE23O5j5IBxX42+iTO3ZDxcAMNc+LHXpLYZEI4IqDn6/o/eA
cQ2rAZQBYNHyMUvOJCMbBaEXO6I2NAcoInmxvxcr/2yBm/B0ZHVjygsxpjE9cOKX
zM2DCdYYSFp0iBowtzQG5Ua0BvLb+wDGp+wiQTII9YhRSEx25MVLDYMXIvFNV2HH
c8h5lOy4YH8DSdL8eorVAsXOl7iCn+kzbsxWesAujG/EkjoKRmmJWiN6DDzn4r+Q
ysvLMD0b124fxsQmA5UFYGEwcXFCUN9F820kNew1AqilD1imO/RShMnT+96AsyOd
5r4yFWYzEbDv0+GvwAwjbbBbaBLAfdaM3oGNJOm7xCsdIpuCozJdLbWpTbf515me
kYVGc1qzip8xqZuh1EE9rBcSjQrC2rr5gJDmhb6geOBMfLrdNpr752w76fpyv8C/
muiucTqnD6xfV+Pym8posWNKBbYnMtrSmGcZkvZORqh5ofqb7/x0qcFoEqRgKjGO
/r6G/3JioKWu+3IBKb8g2go3ypHwBXKlZXnHekGT6nW8V9D4QKF0s/xZBZyK05xZ
KI+/sud6aqwNtExiFw/cmd9D9wWdq7YvB1Sx+Ri5iBM8TWl8m/si7MFjIJw+EXf2
Q28CkxDN4m8yP66ya6aecKSOIJGjjtM+l/o9T2YA8O+bySSsWSK4HOoToRXaYfif
uoD72pT2iCLXMBIJ9B2E3T7e6WsPemzBEJRenOIXrY5c7++gEdBllmD5mcDNCV5W
acAJZZFj7LZzI6TK/YAvZj8Sd9MMsTjFGUjLfSlUndvPDqwD9MG3U1UU6d8dN0UT
H7KRs0oWwGgaW/9KRZS+e2jkvj20YNFntWPJEabzDGbJ791fx9UDsQ6QH2idN4Sc
yU1T+b2H/GVe2+Wziy+CcexPUnBlNkQhb3Ts5Q3pNPaO6xD6h6bTxh57VLRVgBf7
0cLnxuXBPTD1wMZ+F2e1ycTHauYUKISl9fgBJ1l8W1zE1AJ/wXxc/oW0yK0VHGih
+UOxn+1z7EuA+E/ijNJFhgSdvOe9AixdKGWt6pA58aXZnzH+Otd2IxUYxGtLF76K
b07MBq6d8M5rHwO16RF/G3B6FNJLYeU7eqqjAl1clq14piodaa1jChzoVcAP7WwR
humyhPAsMHQKlQOk3gNzvDaGLAJTUAZ5uru8XK3mGkVrZlpWwh26nQyumyfDDAkv
pVWrwpmD96k0oZu3KjeLF0PE3SwSQCJ8LZ62LGvQdFX4WaI4KDO+GNH+1R/Ww239
SKSpP7Ky53kS+EgjqKkghj0OwQywoXMhdhbzow4UyuV9ERdRJQfZ/WJhiYEEAtBd
laQLEFhGHfje3qm8xIOm4CbLZEmIGD3+mXKDpPc7JwfTXhQJNv8DcTARUtaXEN/q
whEUWCPytmaYOGQHVOwKESsxin+DifQJwcYhWxRYuAsMaY2+noMA/hb6nhViOyHm
lgm8iq14ncbXQBupqzk29S25opas6XVUA4aNzy6oX1IrC4JKMt4XZxEUl97nRzze
AJS0u5SHpBO6S/xpTQuCtparr1ZJq9uSbyYz+jPkbNMoh/Vl/WvLHz+KDJbBedPJ
eA1H1tvG0oPId55g/OkQKKeRtWoxzMecoMNm8tD4/hPhOeLaan3Z9qBU8GOfa0Fp
GALX7CDZB8sER4ifKVAy7lWAEJh+6Cd4tHxgBuwfy0G+PEtAkR36Zjaa5jQyLpnx
yWPVbab/Ox1Q06kx4a/90q5DLhVIT/Dx60HpvuZqnoAJHTfxs0K0e9KHLRpMTyuA
T81bcv4Bnl7+/TeAoh8WA0NxvDDieoEn6FOJGM5U2DmhC7+DN9GUsXRSktRvLZk8
ewoDPnhHN4sCZZ2mpskuq77+SmtwozuYD/4JWqFQMcgSUBBsaSqEOA8D4JQWOldQ
kqBLkGIc5hdyGwyxtb3uG+Ir50xDofvID/pRz7VOAGsxE1AMA0Rf6fynE2yryMlb
q6HYZIpWAPQ9lETY7DWLy5k1uLsVn0aIwFq+Vde3Kdm85WnqkcRbn/UfSE13XM8K
+abnyGaMSIhiAVSdHVbGBF3WjCX6RTed/h7ZbVWwIM6+rHIzN7oYvLloJ7r4ZasW
B4gRPUvTBsOIhRGQEtWXYjkj/C96HgKrVRFzCDHmTA+Ud+7LmmDXsJiJiq8WYmG5
CHEpUrh2YSeIIJQPbTLwGIBN3h910bILlVU6rqaoNSsgulgcRCosvqqsd501/yom
+k2E43zbXwOjXtRn9I/0TDIlpGrIPSFSBxl4CdCeC6oCq4j1bMXLsFpOJW6jzdKR
yyuHM6WVHNoTvDg48qPjiD8JpZQvPdak7zSqoqSS94qX4OH2LCVg4rc8Ntm6Ey4z
WLjTEesyH5R+f0p1kNP0Z6DbIr3KZYCLHErga4PDZvI1hPSCaZUT4sA0dwPFL88c
BTRFFo0uHoHRFOI2mFvEyRiUEcWbCdWwDlQKtTKct73R19lfO0ie+5kQ/gFl++i5
e4T/oRbiI5CEx8OGP/N3azuo3EPa8ydWa35WVFQAbXDkr26oDH5DSK9BE+xebd90
DUO0Wi1l+zvjL6ndaomSoKNMj3i/grfnh4hMFvRe5t15zsRDaO0DaJ9QXOE4/gTj
YittwZHHcS/pUSZT86kryJfyDgq7BFBzW8UIWz5R6iXdthH9KW1n+cG+gmYpPcXY
FF6eib2Y42j+CsM4Lo0NiimjAzzD9r4KpnZm9oNXz+xxg7MFugMEEqRkLEVTdQaj
2Y08ebmYSdojyLEgTWiLubMhIxuTsgzlloHcLtVcErmstFd4/UJjE84mdPVnYLzy
/b4WDazKW8NokTJ2mjuuj+SfDY6sIuSDnff/dumPrvsk7SSLca/UEB+zr4iSOixL
cjGjbBaIR1xw377X6iK34ARPfwI4uee1X/AIyR/EXgDsfrUwNcffmGV/2BUxLC9y
HJYbxkRHUwUvjTqbhrQjN9yyCb5RPsxCx5enYy4RPxbQad5qPk2NO01Wpx8SGYRQ
JDP5v78+5EbPyfgblMpsXkbfuDF2Zdjq549W3Pdwx97mn2SiyHz39MUnHYQ/+9r5
nXtWCvex2p2TkfsPBO8rphxtTXaBcpZAx9u9HYrXOmhW6/qIbu58zw5xG2UncDjd
NT/j1V1L8DEixgY3AOw+tI6H979Ijb2t3b9T0fXgFs7lohDvjj3xzRagB/exHUfF
xOKL8GA+0+gZ6Z8ycnY7ETl0wE5jQlta9gC49WuE0hbCIc8xahMkpkAhPLCohwyR
7zvMw5Z5BSTralDy573viJ0O3WMjts9GFu00/D3mw3Ov8h0CtbPpHZvE8ukK+BOR
xrghlGlqWLstl3VuvURVTs6PkRDFABzzJjJNizJckC6xZg6cxA9szL1rrbeJgBLH
6oqHZnGBJdxcXDLCzhQQgS1O7RfMnHy0GZo8+s+CfGGY1arJpOqWKm8YOi0HLi7i
+QJHOIYezXo8hoRttcWViNhHcUIyvVp0ufQxFZevGlPWjMtCSQpOgwAJJann19kl
vXI/YXZP/G6lnD8myNOCvy7sP6JeBW+qs0sS5VId7Il08mXwsTVqL7ben8AEKa/6
nAuuD2QGgI9fxAGgEfLjONUTGT3RoJzHKClcD7FP+vCd6AhNP6PylTaxImPRGGCk
ewTPBkjixzv6iUVOoAjtMP914Kn32LqA5gI0Xe+1osjxD+2ErOIG/Q+b9swhLknV
7MYvvTz1sZPhXA9k8XhHkEazfHWUR3+1uMeqhxKj+0yZNuzgJBg2v7S7dLPZz12F
4zN7kIZVusaR2w4CcxXTWlg98l1scyvz/tmF7MC41mpdUVOomrlbOsXgljYA0wGd
WPKFkKqvG49fsY2mj4KKiZS3bhIJ6pBMFEoPzkUD1LaCPGi5nTdbwPfwXFDDlfOg
m7n3edX2nMGHv4BxsX5iOLvrvdNWGp5S85w6DMy2M8VKXDyZeCeSCZHZ7V+qkoDa
qE4eLQg2GGQt4zoSGD0qmPp656rUgXvFe75mv/dxcJdJ5utVK/QD+wzxuIPSFEsW
Oajx6w3S+r/u2/ht3gLKTVaip+7FcX74jc/gjjmb3p2A6Lt7QQandhf/JV/3HMDg
U7jZmrmaUqUQCBDQCgKxbA6die5758Z1mZHTiKNrS7A1KyI79kjvX3EuNPI5STvf
9Blf/yn5Bj38l6/xCGL50q619xXIBcej+XbFoXSuVY84q5026VPqqDyKwc4pAc/U
b9YyMff6uHqJcuLbuFCGUqvKjYTDKbtopiB/fs8xaOKL4D5Lu3vY1tasblGbiCl4
JQXoWboDGYluWtxuib/wo4jOaSSjbwFGZQxJBZby1dweomOKhnpTZgKZDEDHbzlH
BhZc/xJ7X6Nltx4FJDMn3h+NAfC1JHGvAuOX+3Kx5sKfIvlNkf+8gtUzYlJuGd1n
ZuRGkcY7fiAG+y74saiwkqE20cdpRQZhtnmr3uBeSGiseOOsgVpvxHuD5veQmt9M
pDQQPxwHJa/uXFgwUcbZ6YVcRpyhMCnRIKUtsV7/9d9ELfo2keNcnAsvJb/7nyOz
EGEx1dda4LPLq87cb56lM9XiKDjPY4LEGxmjWE9HMSoffhwsWfB5P9Bl563sDkYl
snUlJxsO3PVFg+KXGB0BUI9ZFnK65YhZjXx1+nH1YkRiZWE9YyS9W4/VOh/XP1my
pN+mzDnR7GqneFqqqgmvm0UCSsj0EhPb5VEvkEzCwY3lucmTVnyKr8ZllkELmmM4
9LgCYq9RHql6yY/kkRXR6WnUm0qN5dEDAQLoBzhVqScrMZK8uNcwiYVSA6tI2ypR
UCUD86ap4f76B/d6hz+YVcCZS+os7WJ3LQoMu4O5wRdV5HuYNV+xLGFJhfPd6N23
s81eMc4BP/vD23aw+li6R2G3PnHgDFbBp/vj772VUGwhkcuZodPon8BjUI91IfRQ
weR/jetgGUvYJbswFjgYNaIT8USWRkqnl0QC81fro+unijFWpLsT/DeXZkGmji7X
IFNCuDVeIjI4Qact3u2XB8c55FuIhM41f3juuO5cezrrB1DmGHb/1wtC7JYMK25i
pNTvPnubgEYpfucmzSTn/Q1HCVrYQK0xJx6+YVXE4dkX2jYDaFx4Yd+zh2iuKdH6
Jy1FXtH6ec/802IUmo10lo89n+GBc/WSHXgD+o0qoIwbdj0a9LVGbsMGeBipyKvH
ThVnlCWOmgTKN8yyVLwjdlSVBOExdSZr4O3WIEVO5FBmz6wJVTc31HaCVF/1vgB8
BnkCoSawC5Rj1HwbN9BxL+F6Pa3nS4+Eiq4IDMYo9fcuHdiPKh9BBQXl9+sXK6O6
1G5garFV9pM8hd0uR3SYzjQUAjxBeUWDnu9BkIwQKih7b0K/g0Lkqrkt10fe7G90
pxoeS0oGfclFH9V1Ei2CCpfU8jc7X/Ifg42G+iKBW4rH/8e8fpyhNAxC7IoZTqTM
+vZ7PkQ5X3GuEA8Lbjy2bhsiFR5DGq3eKYb3uK7msnhSkr3esReAdo9zxTk4jgmJ
TkRSoomJCz1J09AXuVYBODrXjrisj7jqXHQtTv/VePvkYl1YiIFVU7948ImKQsLf
k9xjxnWoY8IxxBoZnorP/mR1mnHo0RRxLp/gk936UU5hSLA00nob1W1tzLUi2uat
OBzXm8/n+bf/XWsp/Nd2otp4kbOuu9Ix7lZ+cMRtGuTDjncJialJjk9esLKCLIfa
7diVntF5y7dVsGHhQBhJcYyhjUHPh6qv5BTtl8VVkcK84AlXU5kTuGyRvO7bceNv
Kpa+CZ/8X8NR4ZMXwl+SKx678WotpKoB/d3iaFL6WO+ADfq/viGv2mvhRz3h05BK
2zMMxsKcBXwJe1P1xDv/GuXgBt6T7ylScasLdTK5SG0f/rJfmSU88zEonxtUXlAn
9eYQwLg1vSKJl0JZLYa2zSxxqVk/yjiEDZtih1UtlsnNKJAQvt8AS5vkVy4vPmOh
OUx8wf/pBesKOY2RsPJFGjgnyFWUm+BCDaQwYexwYIdcIBmKc4ViIRomuw/STJoA
OJNBGgn0TJVc2HBVVjVzEW7vHK6FzToM6vtGiS7y7XQXnZ5ctLpV+XETeZPFxW8O
unZtR/T9ekBG5CLp3ToF18A04+aIgf29WpyPLXnjmQHvDPei3p2Qa235+lxOvtKh
QKcXKSyGthfbI+fSQaS8T3LB+4d/nPgyRhhLb1xHEAu1u6Mofo988mEX4S2K9nvd
dE4P2FDZUnqyJROzfctfOrI0k43udXgmk3s43F7KElLiysrlZHP3kqpH/eWlbAxq
ZNPBtLaRgxoX0vcxnkIcf+UREVG+diNk99iTXGs5AHMVvy6KTbUg56Io3aDWhayh
jj80zAA0UJHeJd3NAGKizjXzbPOTzfWtgHezrAlmuqm86aJOW1XiExR5JvhOljGU
z1pnhOe9dOhgCidRPS7gXzEePaPcZOV1Cq6ytedLv3HhlcsKZyI/BRmsr9X/1T5v
jElpBnO1w8UStOMMPX5ZdCpKQGDMg97/w94Dwzs4F/hFLFNYuVZptsS3rHHAUbm5
uxQRjGT5m90cc/QbpCnAkXCh0r3IRBeWRMSB9UD2bSTlW0OCMw+YCprwncK5wdLm
bdy+SoDUXwj4imGswJTyXIpb7rnN7GBSjb6TPzpTLIVCydnf2+uTUBeSek5FVnaC
ANFoJPPPoVOZEcJlGUxs6SjDZo2JEDwdpDCez9Acm9KHrC+wgHP9a8aWq0WOjV7q
xTBQ28UHykEUePEygQEV1RD3X54+ajEAsBUZrPg8rE770KbQUubB/C7hyH9/QDrw
sqETfIAOETSIwx8tVLqDUFpIR+JWvpBYs/eBUnlXPxsCLYQhZ1V6Ff34y0OpLuCN
e4f7XHxMQkDNi2coEtWLK2T8asoWMSynxX9ikksPOeHyhdlw20WlyRpmRUa58stm
CpY9XsfUcbA0T8BjZrXV19IpVaXDuQrmzsDwc8gn3r6GvRfns4avY1nabZhXwHnO
kxZCeoYMRvifrpR/Wv1zf9lmAov+e16IcFjFDfPP22CXpItQgXQH71dUvwvsEUWH
C59cGN2ms7qiuojRIXTzMPtEg4ov4I9/XgaSb8NdFfUo/mIs26hHJw1stdiI63ca
JGvd1AXCdBjzRRhUU5+Rq1PvzGej4I4Q1h3JtvKXnazjyiiEMV03uvNIuxTc3VWd
1in8+QJKACwWJdnnqyaWUZUyiO78Nq/shOQs1U2ewsHHr3+ZDQOx+AV7NlOQGKaA
uxD1+VYZHzPZ/KdPLT+jaeCCV6tvOR5gyOoGQYjg5LBE4EfANfy7e91O1H5mNnj1
ctZ2OZA3drglLBp/H+sC0ieqYlgQYYK4+wld9ZQg+7P603qg6T2QzdnJjS1OoKlx
7Aww3n7qbsoe/TFoq8m2/KfBlYaLOHtQAw1MJyhWbBiA0wmPJvxCxTH13ZVRdGND
oLZGiaI/Ns+9mC7/G0o+9WNHk8AGnFV7+v1z6/NeHAVKAro83KWUfHLgpiB5CLHV
9fLINVOjP1KVM8Xh/AnQJJE7jQtcMB+XGhT9xe1Q0gnm4sRcBtBAJDj2bKA+XUOl
lDtrS7gi2zthGemjqM8p+t8QO8XQoBQfuK6HUmPXCkY40KvCLkkXBCEhINICH4/I
RpCxPvP+aHI7qj3aiyAeP7DKDHuHmTNbaYxZcQATUuLz2Azub01J9GBS6oIlugv1
bNB+DFE+9qm3UNv8HLGgLzrzGoSw5qrpE7PSKEnID6VeWTHYY/p1WQcyNITmYXyx
e9BIwsJY4kbXPEWaBqfTfrCuCPS4fzsUcCnp5L4DvvwgeaWFwLsVfN8BXaC0f+G0
Of5ytkjNWLmgbIu0YPh3MDvWJmplkuyUtQvUMZsxgSw1Bekayaw7wnmc27gCTUWE
L6ixzsjGWr3jgV9o6u8MM6JkB1imEon5WpzPh5Stjf0BQFwTYUzaiy48TNAiw5Xu
PhjiP1EdEHdZgNRSf1k1Zowm9OaL8Our1GC1iKCmTmb2zO/xuK2uyN00RpGfWmeQ
dAhS33GQLNX4kpqPyxHkkYhxXdfxNjmdqApjTD4/Xeq+n7WvxI+re9VVhQXTHXAN
P32wRFWlqzp61auWsyMwy702+F8YtKzYwZdQZKGRc6V3VJqY1VvVZncZlEA9ijtD
aTf4y5PM819UVpxWmY3cCv7xdbz8nowyLtxx4dL2qDU7vUVUhWG0Swl2YtanFvZU
nOCpV3EKmHyaQoY+anKqsi0MHaIZuj49vs/a1zXWqY+n+TrW4ydFdYDo7hg5mWbC
NMxdfG4af/XJgoYk8P5SeyMP/QZzkivDROOp8WOEqixVuEY+Zhd/R0CwP3lqcj9h
1suUotSyvWmDmsAss1heP6KKn5HtkXW5XsNCOgbz+Syr94TZGYVvqrhhH2FcRkvi
xleD/LAwQK5QHLIHxXEDrK5aHgTQu1qWsMQF2sx1XQOESgLkcIQiHoQBuOCwNkGJ
epXC5uRsVMkdbMju3k5SzpUinVAqHNy7mhgfTkQIBqDMyY9HzrtOD8Y1tc2qXjr5
NYF/40BtqsHsViXzxSah7c8d0FGscPYgiAxBItSbHgeQD1fa95iy+0so2bbee/7w
ye50P0xTkZStKwuPbz5vc5JDIO8Lk4WbkfscsUGHTj3YKUrONCB6fMiHHqiGNMoh
iW4b1NeIjnm2RqmQVhevfQDAHSsCzgElgk6qsF7ZhAeaP25u89QF0CArszRP0CBF
+5NfiFHnGm1yL9Et0OYEFdstnScJ87rC2I13uxfdFcV48K+bfCMXJTuyoDzCY+2a
8c88GoG354bLoholy92b1Ot64/GsUjq/1SQCf2Zdpjcag6ewSyetqX8OVLPwYRmG
2ewa4I5t3uKIPOpHb8E72QuEjwtes8oj0Ok+nsBgy3C/TLz5xxfAwrvgRayVjYQx
YQVQNYUpw4a7IodMvE1jnmFCO0wOjx3r/sZGNzuWoV1ON31NPjjXwy9kk8xvL/jt
AlbqXSQvqj2tEsSvAht6gEpEgpheKQ49/nUY7kW+sBGvfMMumi9FVSfFN238sAMX
fvI1Ce97kvoU0LWxMrWTVtqPT/pzG5uALCcgTNJsBuYMmJBwVJE8HAMPmIq1V2Py
F0LvXkGbs9741HCFKaSRdIDCJp8o0DDa9WWZFuJTWDVln37mczeZqA4bSBKihmDR
/tLDdbDPyctYntzHx29bcYPIg2Nq2hqbW+RRXNxcuCY1SSWLYxEVcljtJY5EHxJ+
GgqCoyYCH3WO1/4KBjuiViZSNLak87V6GpV8UN5godUwQiOUVaF1hN+exhuSn5H9
cIB5ODgiL/lUN3+CL8gvtKpnnYhF9eGaVlGgSCEijAmeDBUaR97apb4enYKdbD/I
MSUYW1iXw/gpGVo8QOrtHcIwGr3QdQwWnpQ0PIzFgFVnBbppvMV2qr4fIGkijq09
MbPK1o5vtz5eZHlW3++CKYr6MBbckuBgdo53rKsjElTivTCn8Tf8d5blGLX4KY7t
JU/diobBEqM+LLzLEQpBx7t0i5PV9TUMh+U1eDXKlJLcxt9awrhaM3QTbnDneFsB
IXjVV8bDMyuyDC3AH85kHnW+/UvxDz7af5w1uW/QSWpiV+0gQgmbeIimpTzjpUxi
TB/cXGeh6r9Jd/iZlmmdDN7419jUn0/1GtWQUeQ1aPS9RbuVXRkemZTmeCxbGYUp
k9LqbbMx8iQmIgYIezZpYeKtjuX7t5FpeIYgtc1I/1KcjWLQ5pMDFKFC3bqTh4do
dAQZoBqiBa/IRsVVSYZufyXrCCBF/grydjYesQ5d98me6lF9Ob2Uwy5nGUlQHs9S
90Alkz+2tloKrXk1H5pFKPbhdPk2bq52p3jNcSFX6h7kAdQmHJ4BRgmeqD/nQ9ZK
J3yancTPiW7BrXLcldF+QmCinVZe6i66e44X8issRkaYSeNFGS+blt4M//Xp7Z8o
pB9zN2h0FvOK3cmLhLcgowGeQBqsuve4J3VqrqfaC4286pjpC63hdWfqDz5Hocz7
9+BcQBATxCNY1et50FKQ+I9zULq2zn8KW3kmXI9lg5wPwyEZpsHetNgQkBAqjLqE
3VLdmg0O+T5t4TccIa6xCwPF9cPaeoy6kxQboeugtozWpReN2huPWMY8TDVvVvx/
wDmK63LyLUd0xfTaCRRsBcL5q2HoUsf63CyRvVrAHGKrG+ev2hcm6NOeAwcj/Ozs
+s5anWH0SpTmZnmKsVG0R4Q0arHEgTyH8oCYbCoTcI71USXBHsBO1RbVhqfb3M2E
3yphg6aHcLfG4yM2dGF8OYGjRYyKaAUCLEcjigeC5/2KA0oNIyM7JMCP8rLxYpAk
w5PGHLUWADRHOXf231GsRo/dZifgQ0r7IiTWiGLaLhjENNwmcIeQ3RejA4NrEF5c
hrJ5joyVzTj0sy0ntBvAv9gSPIZzFTJ+gLgo/R2ejCX1v+FojhDT3DXYAbINw6VF
lI8VfHC8JZ8Axvy5SNOkOZuENbrZpaDil0Ug2GFGWuPlFCYIWhN0oC8dPjxH9DOE
+9ubkg3c4T6yRa7luiP6lInvgHI3bIbv5gRvRbRLB0FZS9CEWjSDtijwtz12dKrH
oQBz8x/9q8wZhDsKbfSNESJeLq48Bq3XBpFc2npGlLszehOIMr7HXVmIuczMX8Vs
DGP+CoGqZ3Iq2oHpVBw31ofd9z5AU7W5QXiV0fHeDfoieF6s89grWYeWq7eJzEI1
xJrTTsVR/JfDUfMwgRjJ5uaTCMKMtOIG6PKVfbf4u/soqgNMUZhcfDNc6J2jWkgE
QtBVGdOHldTgkOvyTxfGRdsL7oXAvERJZiWhL4JQW4RYiJu3vyJ4z7jZWU1aW1Jq
4NW/O+YqCoD80YaBP57wOeSkSWOugwB/WdMEg8JKZnsZ6MiYq927lP4GtT7QGno5
S8bV/CDXXypi41KTfsNdfh51/b4gK06ETb/EdK4RNHfYbGdSK+igIJQx0bPT2k7n
0mHiiiWebJ7K1OSG4i9xSUNg1re9Sj/6kPlF7hQiNP8Ll21JkYgMhoFp3Xo6HM7d
yexKm6Zx7dQKIa90yiTJ7IuWQz6398NrS/1Ye0MCbsnOkyDlk44FlmJq61Yzm5tI
D7wqOJMu3XlKwOR6Z8MqD0q9rBrVwW/ey1O1owexp3SOcwVH+LVL+W0Pj4yTjPBz
U+2v1vAD+BHgSDFC1mS5HIB5aJzcaxBYhxpkU/7edZWa1VQGDsY3g7ivrExpZJwn
gy+e+TgmJYeJ2bOYjwBKV16koZOMSg4oRoH/9OeCgWDr4qC5MIQ3IHF1LZZEwFKP
fpdAJFP9NQhJTW5k70KGB4gVjFTVjuqL9JOng4ArUaJ4uKsWnJtfpBsl1qtDd8eh
0CX+Dw4U3t+qHc8xQ8nMOvXglGPIE3K8qvvhe6zxmwmQGTqA+jvEA6YXfuNANCl6
Cat7UoOPMKXnCpLFHbj/mn+w0doXsPzR1mwLfK+lqVKr9zdejfuLrsEhtJGadSm2
MoUevAKWRa0lc3qexawBZKOJfzVF0gxCw/CdpP9PaZGLbMcD3mIhmVO2j2mnEoBw
PwGiAV9QljLkfijo+vMr0cUU38pPdy1csLzZYDpxtlaVncozLXtrIc9qOS8AJQFF
2HhukUCIlWUIFAICjvt0T1TN3ST32PkAEKDVWXoO/NBvkdSqsU8cqfizshYQ5szU
H71AMJE6SYK/9t08puoD3+Ha+iPCsAA8rkc4h5O3mSJVsp5oXmPVRgkD4ZecdjyN
uYbjB8uFNLzmD/p/yXQuZJ1E29GCdUSGyvqZGPYiN+kKKPHM3ywiQxzEwF0tF5YI
fuuK+9KeEA4QI5K845rCVjXl861v3IH9GVGmnM2fv+dc+7bR4Ve87daq2D6dpzUw
s4c9ib8o6tFUx7wC6ymU5jQ/sbTJBMIOGuk1t6riN1LIXk6ryfAevNHauvzK3mj4
BmQb+Mah/RYFiHGeaqKiqxfy3BQIg1A6f6DWpjPEQ8l1wk3g18sZ2gXU++Lq7wgi
PhtAy8MimSMeAMIgu66Q0KY2C8SIJ/mNo8iZHNe19qZzscclmreAm3f6/zaKCFDe
pNM5NHZCWm25B3XGHzHWhJZm47cFeieATy22gclgtDjjVsT5bO+6vFkpsvhyA7WQ
6jZ2ChMhwXxSQfnKh0zmY4sfQse5lCddpg6BE5/tFQ2bRm3Ki/EL0sbschblZtg7
oGu+Lc8jjIoS/kfZrH9zCdmqsGfgyzeLjma/xLjnyy5KoWhHV0mpi7pMeL67TLkE
k5u8X6jZ54Th+06xSrZcq1E5Qn32t61xtsXhiU56q/gsyhtwrMgrPVQPFXopver4
rbVDTTMZoDLAPtwiKMUucxeDi7ju0c322vnaBi9xYYBwCqooLUL7cC2y4gAfbgwC
/oM+6of2M+ImVfsi7GM04OzHw4eWgViYYtYbBfGfseMtNNor8a+skFGgvZnldJDF
6y0riNoENwQKb55G1/sCbfa/mI9ggbqRkZrmS0d0QhCkrO3AY5cvC82Ki3zkdOo8
3kV1Ofui2zgCUq8YKfBrnHK/AIUVYYMRuvaUF0ER03uIJie29f2rwV0fDQ0JGPxZ
vg1icXpA39eXfcU7x6NfaJeG+lc3XwbHVaG2ubKyovh4sH/ugXTJwjh2l2bm5o44
agavLwsV85taAea223LOPkxrIvYZq2dxQDAS3J32i1xgrT5h2Y4r2ULkgD1wmhrf
chWlQkoHFrpmjk01TiZvZHaiA6lYPF6HNfGRFg/aTEOipq1txuYHIf/fxbOl51IX
sw9fBCaByxPTFBySx7Qg0e//V8uFBL/Ay5+Lk2mgzIRpqyYycwRkHeAps12Yl3Jp
QkjhBFgGlncKRJgvjTuEmu1YZycZogxKW61cK4QTU9ioJgtMJz3j3MEJDlpvpePs
EGE1l+e9uGJXCVH0CDCjQVFVJJ5PxkUxVVP0rcZmNY/eW2TqwQ9OdiVBIDWdLrHX
ZLMMzg5RFgPGzKGM1VzUJcXq5n7/1gLoMxegGjp99HyYa6ygc/0Q2OZgFaU1rihK
kWKTn9fYBzEBs5GaO61DxwDsS8ZlqEUkx4yAl6lM43cT9ZKVLXQhhIIm9Fm/K8vs
oq5YTXOomXl2aAyXISUqlyMspKLOUxanpP6wToybjymUIlZ/Rn4IRaKGU+MbT/xu
PDfw5tDZk1ZGrn+d1x1+qTosrYKvmv39aOujJEjPFnQxwBo5Q5CZ6/4qKB8ekuss
6pvU9YSp2dZGtrMdgPObXHuY0hYEQynCF1lKqmA0Imr4dcXFX9HCph611oS1sD1U
cziHQGJ80MuLHMCBN567u39Xfpcg+jgyGuKWYJxvSH4bxlJqfTQMKiZZG9xT3Wog
mmCaz4Afcw6iASmtGeoyhS/tcHwrMrEruVkN64//dxaDbf4ArOrCKcA5aVRua+VY
oZMf66NTrxpNQcQhPIswLDXGunYioT2bjObbJ9ma4ofNfAuPscMsdf3+n4fGnsdo
D3AdzS9A5Cmtvla6k1G5Fh78Wam+NwXQTqNr/z0ElDdeiYr8LM8O2UZDsBR6jCx/
qLT9iX8zjtvL4ZMcy6IYPk5s3M6HIXcmEDtLW2C4gm1GFXctSluZ0WAXbpiIHGvW
eQjC4UDZoc9TbbuVYuog3FVGoggl3YaiM+G4jaqOEnpklet1SKkv0zn/V29sDqQn
KIyz/rfBGC5Xqlo7wdY2V86BwjC9j0mNA0WFMTCZDCEvzNJ1xpkhUtyb1I0cpWEC
RQ/cStT/2TdyaQl8Y7b4qTCCQy6ksHVI6beZuKypwUy2ZQiiuQCsAdnPUwmn82Xj
PUatBMcutYNfZ1FB4lXrnQ7pf6S34Ib9KXUGj3RHubWps4wO7p47B5v8gALyi1BI
0HQqcoAyVXOqm4lx5OZeOfzjHoymCcO2pbYG0FrnVQpB++QmdRMzrw+Nsy+e3BE0
j3eHMt89i0kHDSDNaOcaHawfdGdHdkWmXC7mdQxivhuoum6rgWt15Yt4Vf7S7p3t
4yPWcbLKBWugjrUOoS/B2OQBAarDYFqWsQHfJuPrTx4l4HrsOikmmbSZYDgXwzT1
dn0kGfmfPw8wUZmFcxxdiGp8VPaBamK/3s5v7KFdT6nduSdeYjicc0WMrssdJIOj
N75iw4wiGagtujrAQcy03XsHH8665V1/HVrOKsNplZiVE+p3sX/cBDt7HhGpkFM2
J7iRzUkVwUrzMgopLrvf6/9eukXz+YgPVFzoVDuns2YDkQZf4QeRa4uk52tuNCvW
mOWwgm1B0rkh292h2b9p7E0RsxuCB//F7+GQJMevc21FBty+H/WSDYFzVqiV2RRd
k7PyDSe/Iumh/TlUFlxaAA==
`pragma protect end_protected
