// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CIofI//9UAdBExUwydX20TDB5cELwT+KXO6RukfM/+bnjsiBixIyXZYwBNmot+E3aEjgOB+ELceG
5bC47luV4twFZoTWRmCKTWjBO1Sg8iUKzSDuhP/dQ6cSZsBShh84ucxSs0GBmkO3ZHLs8dxpTVGL
BvuG+TY++mSDz1PDIfFcZn5mlVE0g5x6t5s8sWKyGP+iU091PHx+31Jte65icVoCiTeLlrUvhSpT
SgBJ0lTMlH9PvHTnw+v/CNCsMLq7tBXoAyZPKplYrYbzo+09ESQ6iSK0YS77EJnxHPdE0viIMBSk
QwRiQJnk2optYIL2QHz/26yewxbhrgVNRY3H7A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14000)
dWuV1dMpFLbaxf9yPz+8nl2ZuyxfqvI0ouhboJ99Nx3EXmFRACljHKWk9VF0VFH6oNOk9zd+r8Tg
qHjpqUN+VrWqTVD7H0kKVNNSyCVIwlDpPrEanQ/9dDgc3M7jRskot7tq+BaN7zy/LC1XMSu9D0If
p3ZIiysvmAbEYmre+tKgdVm4n90x2nImwR0Q+n6QbIxMpaO+K8DSAUfR/ByykqUlab8n1AjCun63
xhzZtfasO26HzcHta5wBNDQX6pygWwWSgQSM1JZsRSuAhYZx0ImJ5Xuv1aDMDl/V7ocZQif9F1Wx
CJ/G6N5mlzQF9CoJUopAg9BqTTGJMsp03TQ5VKu81/rBZnEgvkqytyZHuRzn8lksR6tvrvTy+iYl
zXrCGcnRHisTSKSvp9HIEzqtqEM2L6gfZzwz96fahA/Pt0Kk9wuVMSVeOPedEMhYIiYhfawXwzS7
1u2iA6/nmMenRa34elAJyUw6WnffSb5WJIoIiio8ymSD/JLdJDsS+pJXsDMMj51VDCqTmRDeO18F
yMkbsCq+GfNKGbQMWZY54bV3tguSHm8+37ZyYM0HlDeCOMNNTxd54qOr6Xd4ROW4lxQYagaPdSb7
HF1DC8XN77g+r9idNFi8CBCGjiErdtC6HW67fGoudwXvRdExQD1wJ8JDDgWCvXvlajwMZR7TKzEz
BzPaFwrhASBa2xvw9cMwTf2pCfhEoVuNwWERSUrVTNrHhK1yAZeY1oPCNyLKv5kGaJ7O0deqPeMH
fU+0jBNCO5KXTKot9RPjCVwtvGonzjzUqwxdhHQ3wzpUw/iEyPxZL5S9Qc/R7N9RQyK4H/LEt2Gi
p/CTxY9fqssyFg4eHmQzcSkjsVmWHTAQ/575/kIx1mrgRvwslh/PiOSK7hTdMSddJ6EEbkA9nCsX
indm7n7PzTFzThUPGXpwYo2dNdZKI59eZ2MAEQapcdOhMTedMk+oX1ACIw7lgfNpkjolJicOeI0+
XIvnpxtdoF+DY2cr6/Qq3e4oUB4UAjEs76INcu9l68xd9Fd8RnzMahQ9Ws1sTdyjPAVXBU67PKNL
1vwPmH8xtNlxhJFblLzmS1GNewd4AFysXYX18HwgebVww1S4o7LohSAzOP6IolT73XK0UB3XrZ4Q
/+77f0hCmn7r3iCCIEt2aHhYGmM8oMyPk6ydRAHK7k3hmb1dt/EWbROKIbCeK5oRpHkVSbJ63rvn
P+URVeMgp/XNmsP8EUcgm9kO+MTgc9hGBOjMqZHGUYKwtoziThjmydyL0y0/SSgwmOd24j6jv9/W
q39QB+/0oj6w62m8foaSoR4yNwJXIw1hY4pG78crk+pyyfekbRc0yivz3u4wACelk35MJQ/CVPX2
EYsPK8zddimPdCwJOzXyH+iW91tiOzPAKdmBoxT2ZwF9ST240a2S8WLE6aLeEvcaen6bR5lAtUI7
liA4wNs62mUy1S4PF+e/+pu8O63imnCb72Nqw9Eth8pO1hjFQfIO9tMnYixlEvHNjQ6kQZInUIkp
Iea5KCQmAjC4zEE4yBUoQrcgD/PdMYY6WHF2c4TPe8LoQjto30aELke72BK3hV/O7ir3LYrS9ahz
IHzG26XrSDlLR8ask28dETsl42ET5MWxjPehSYnB/RAwVviOS/xTI7fBqYEZgkqwPGAJCp0EuT+8
vrTC8SNAcnP9FQ+E4ElSRZc2QNW74ENGc0Y8wHOaCxAbtjtTA8YmktdrXqbudQ3IEqgfZlHt1X15
xP2obzzYlXeTuDXsUoQm8magNjDXczVyFBHYUKOlW4s4IIt1DPzxiI4zdBmLFO9p4OBczZaGweEW
JXwaDakAq8CLhrJe4pPaZAovh1v2+yObNLs0aPI/8MseZkGXhKTBdmhj6EOUzZDriTWre50Mh8iU
pi7oXzEgCg192WTSPPbiwXaBL+s7RvaBsVGrR/cbr8dlWUyQV1Hp1OvW2/lNgdl/GlwOUj1hn1mP
zWN/MR4QLpYR/8O9WUpumKHi3OMyvzJCIWFARyDcJh8Mp30w8lnYMTBFUgxi4SyKpIl6hyw/tZYS
CpWmjV4VPsjZJR69Hu2w5Byj9OH7YM7XWdAjtNnT7tLgW6t4kO2JD2WkGCjjfQvj9WU9MhldScTi
YM0ewPBxhkKt97QVAiQ45o+3RXSIKHZ6afV2YICItMgRGnsM7vDxoz/8/S35bBYxjv/aiPknbU2W
C4J20FcR3/mt+iN6pVIo1Ek8p9pM70hGNraZcds0zqbF/GxAO6FglD42D6nLPWAR+tox4Yvi89Lm
9LblXPQIafzHhr7Rw4sCHxJe6pQou7KeYb//bIJk23d9/Y0MbeQ1GFW6h4bmHhQQVrVkGZ70Hpix
SAGGnUMW5Z1N12KhNCBEnA6M3w7cY1tmVMBkTE8NAy+FWpmmZ5LvZiuWlqFR3/gulM/hHJMmswZI
mG2xJC343wF+yKaj9qPudlVdHi56jppzqd+fAQkc3W+00tfKUPyzoqJOrTUZcxJJU/jRUIPVZnoE
NM6Hmlq3Ba6VPaCmC4R9r40XkRvQPO/XAJNRxJAWOgm/C+U9O42GRHrfGqW2UfrhcgP1jrJVi6OQ
PdYPqUQQpnViRKv8rAD5KO5NHNhdn6icLjx7VPJ/EVvuANppU4HiaQ6eGo9aGXFgeasVhKEHA8hf
1zXCIAxnREEbstVlLPUTdLroQHe7x/2pSp9Wq1MTJz6kaThC7Vtjodupr22Bj3EhY0mJubXRicg3
X5AyboT8iVFrI6YtgT4/BCtcR0woqP6OvTlmB0UZweCFKHAWE4Y8h6Rbt9J2DVOchHA4g9MMGJfn
YK6E7iiyyQ1Pddho8tH8fc8FBP8bKSMGGPkSasAjP1BMicFrqnmUuHTJs8ID6urP0L1i1mnB4h5C
J0aHiUkv2J7eL/6ZoQUzx1xwHjeBgTEncsO9tWXGjKDkDn2I91v5o/hSfw6QTqEVUZNgy1uck5iS
b4T3a57v/mjAxtUNUmsxeRGL/gv96p4DCNOPGwlrhSmEWdZTD+LjofKOqwalxSibs6LC9MZr1hEW
MWBSRTKclfeiYkM/rnIVO2HG9Bl+0RAc+D1aTewE23KqB2t35rHyTqrcMyPGHsLJa99Gle3u48NI
ojQmWqmKjzJmmvC8POMZeFA3FMlf4EqJHgR6szyfEJTuURSKFTuVlKd/PGu0SYFNg38ZJWKYhfSc
eMRjY0C6Bwo1BEQdS2PWv4U5ZlJTs/KdyS7xzFXL5VsL4Kj9ortIABIqqvn+0k2iE7L6OhBYJd3c
np4m9lRdOI2t/hYLC3Nge/CTPkXxWGT0wCc2fs2/hysRqZ5ztqHWuwcIk0RH1LTpdY+NJlRCNZfG
ClJrNxL+rOh/xq6fSJTq3nP/tTQz+74VsIt0LUXDZKfXKWV+d1gfwNCifUKdfXnt0owY0AHNC5V7
igCV/sb0og0i5YI9k/f2+oeFUjhGDbCjdudT01ggARD/JU36QdD2mFG+wlB3rrmeIcfoSvuckZeo
FS421l5z0uSxohrExpyFSbRYqIiRLn84Z1UbqmzPnsS6P+mqB22gWRiQ0TcXcKF/YxtNe6HSwLzM
mV180n2vAB94cv/0wKUmNrXkaWV+9N2umYKm41mMeffc2n1VC28hwAvj4htkx+Pgdqlccr2iR8PA
42KQapFTFSRjK2buvyy7guZF1UGV6VvraHy+HqlYatlXalqE00ePB40+bcwVuHyUpQvrPBa51NrC
d1qLJTtTJafdDv0wMrw9FJrePFy2jin+Z4DVMRTXAbV12N0ItTjfkLPRoAncYe30RytJu5ObG239
eloQhUYFzV01+rCiKUinkbeKgy0uP8YMDHg/TrCO6xQy8LWowEKukQ6b3x6Cb62q/mCOa1HtY2Mn
xXmq/BamkTpXh/vw3oGm8dd6hUEJ6bNrKCRLIc5IWMBxj80BUm09AphpQTdFH+vumJKRS432LRqx
W5Z+jnci1MxYv1jQ54bEu7r22QRUEB8Dxq5V7ebzUdP5Oxg8RamI4rBaCJ0eGI0uqsPOvxEW5G6l
T8CF6G7SLbFLbmE0D5pBFP03hHFzdOBhovEO8i+B//Mwm3srU0z4Kh1DGrC1+boyhaIUOQryziSk
VGwDsTYHPcd+CmkQ6fi0mX/2ibgUVYJrWJP7iTBLg6qTzIkKFpYb2aEyIJX9MHge1z1TZtJOu3A5
qcXHUkMWN2y1uWCFvmj3lyshVmFPkaEfGm+Xk6/JsS1PR3qOn7kToGatlCD0priwLHnIuguTvkwg
6nXMhTtpUI29hyZuUf2XWL9/83BbG6bLuRnmJwQ93nl08w8lOjrYwOMbr0CBuxf8ttQ8EMr2bAkO
Oc9w0e3FHc0zTrrGull0g66dt3HfJxy14XoTaZgcZhuVfpE9hY0MUcX5zX9PZocAAP0EuiElyucH
02j0xfZyLHPXa9ecRhO21K1iMCMLdFFWZxjpZucsM2uMjlHHOrSdIoRgbYjx5WhgLjQIlY5sWrzy
/5G3Nozb1kNSe09CDDuc0B13EaHABD+68a6OpLxp8tOa1U1yoHJJl+7vThX8/wHT5sE9Do/MUrTy
YiJm5lnkHtYCy4bEn36l0R5agWXtK2dbsj1wRSnYJVURoZUrKzAYxmPLH01asoNDSbcFOsEALFAp
rF803nNtWdS9+AUuKUuXK0VPT4kNnGHx+YwJ0rV4FQjj4YHDF5h0dsN47NOxrnAgyt1mFuyeMR3Y
n9e30KpS3Gc0otVTv5M5nu0PqkNnEhV9YZXkRzL53v9wgFr5fZcfAEg6wzxcXL5bPvmV0Awi8zn1
mu4lNIs3HFSwgGBkm5WK69ZFywZ1pr1OyZS56ZwO3a29qOItYMWp0wElOe6HP86FAasKQLCyrTFf
i3mAJ1JiUx08jk/C6dxBrCDaBNlOEObaMElO3EnDoY2R+BTpA0Gg198JQur5jHPQCAuJ14cM9oiJ
xdjg1J7OnnxEk9ENm3pbNciulPjZZSPn5NQPVV8xq4XlwH9Vv0N8oeUknVQ2KURpCn+3GAvTiABT
H7110p2iWT8aLZSSj6IaZTDm2d2GP+L4Kykkd724ffWMbugugjih78MFrNjmau6eX46t0zMgbBCN
9hSplr4hWSR2yFsloYdoezCyrQqVZ58Zl8fF7Zb5nCMiIL2zK3HHcUtGo9YH7O65AYwSk9dbCG88
TQJvQMgi+3QKG9Fex4HMWnTPsb3dSngmR94H0KCwpvwD/LTREYz6316QXk8Wlusx29Jyt/N6k2lf
h/xw+GH8IWx9LJXVdLwSZNvXZEV1AlKcBU7DjOinrVwMDxibijZhatRAZeeHak11rFR2bU+oJPyI
iSzTak0M8YOwCoW8vrzzm6rykxju6LX4iUGqPAkNVoYQupRZiD+iiQ5IFRbC1gs3i9wko2B3r7jk
yN7UwX4E0/ommis7FzgXUFKieRq2p3ptJt1sTlB6chdjrrcFHzernDpRRFYdLcaq+SN4li7zWJL/
54nIsarAeXxjr9MPW59Zbtg6N6enUyhei7PzSEF3Olt8waN4M1MWLLhybmRaIjFLwv2e946ota3u
aNgMuTD/Gqtq513M4Xcfvk/yk5zYxfzfEzAIV8m0vJwVANBPxTfjT1SbpqLx7VM7k/N9Og6bSlXJ
xS3qqhazTLVbBfE52FBlonEpxX1SYdhII4XHw38oVVOb7ttHz/OPZKbwvyns1T/4jMlTEfK865Dm
XCHF4SXpamASIyiP0S1uQQYAszLz601IHKTmM637Tr+3WdPMv4QRmN9Mu80z0jmlldIBpKvtTpNr
Hta6JoFetkyIlIF43szBAK8XkeT9ezanH9GMCf+4FKu9XdmxC8GtiaBxOqxRbaXRi/RRdjvakgDl
qqyuUoglYOiNsOsougtT9NJEKtN3OIQrIEEeAxu4zfMyjHjG6ZRAGibRxehaE4uokFr/Z/SodSFJ
4lWsO2vfFS8UFeZA02RdhBFH4ABgoLmCno+Ct74bCY0JvpjwoFVa0ypleH/CPmldjTnsazsHpM2y
h9IycAHKwW0unABtT4LJi6xvo0VSsOsT5CI/jvKyus/umtuuOOs0zdNZtXh+2w0bj+AFdUv7z9oP
zpuMOrVzRG+RiRKdwb2pfrt58ooO7knGJVsDpjrFV+jWWPKK4PAx9gxb6Hr9tMECzpBYOEegvDkS
1r6jXAS8xE9toacdZTCUWh6ofCraZaBNjieuNcNURqKJXUZjf6GMZj6aNnYU6dTj/1fsNT/SfdHh
+ZvJG227RPqA6rCM3wPO+UzAHf7E+BPuaPFmkmHr7252VxlnDVdEeyVyK9JFnWEXUOIFcuJHIqMr
hX49n7+9mYt2Gn5UQ82xhfZf2Tkij0PrJhA9EJ9d5u+Mr3LgY4IJjMQVfilirYVIyb0oQaLRvqIz
6ae2CYqvMtJu8se/LKXGp3wscoEILtxvn0WSFM010QV2tTdVomPMkssHW1yvkPVukATVEETF/E7f
80vn3GHp0qQ+zZOBehgNd1Fev78ja56+N4mKulQD/Cl0hzKk//BBIAEJCDxszqZVzJqPjtF86WCB
RMUflKr7aMpJc1om+MWVvB3u9rjnVYzsOdmgHByFETStPQ4Wj/u4Fw7H08jnDSdiVbth7mB6mqLT
4yCVNC0XjFcDkIP77Oyf07vFOEDACeOtMzk1o5cOEXmW2fZQx9JLeXzKIDiUHZrVTw8VASnGCnUI
hRV5FxI3H5+waaQJx+J1sFZiBZz1HgPAnJoNtiZaYXY5uvvVkV0WJ9CF45VUhUCpmVfTvk+GW2sw
Hod1uKWvh28FAXdhncG9qcFoYqkUtxfZvwp/7kQJnHAv3mmBqVgEsZbjA7kFPF1S8UkqTxrxNO1m
bQdNvvEkppQjNq/5VPwVXZw8t3va7hDoSZEwbytA2uIpl03dO6AyCc6GBntvnXXjS8fgTFcWuSGL
z5t/k5Q1bguhxO9TuxxCwMwo5zDtyVLPBG5tExCGsnaTMud0r0FtwX8F8fCitPgyWnDTLPcMtip/
dz2Pc8guqjBRooMsKBqKhLKnojXeKHZ8iRF4h8XQ1KAgCCpqgREhIUGnfsCXV0hEdgMFWjNDATJV
K7Yc9QMUzB6u964tBDVHRH0SgPjzXnbemApvwlTP47Mo1jUGBjAqdnC+IZuwJOvcCgJO8x282o5/
eAE1qfyGtKjZtS/Q89ggXsJ/i1u6DP54kInV/76JfN2iPd6slAkSJZ/233ldjlMM6bMINrSOR66w
WevBNGls51eR+GtC97I8vHEPQUrBAR+2yKMiayfSxe0vjf6exAR71BaN2OLaFMtTqK0rubOu2rd3
4dIbV8UiqRMxwnramV+f9doyWkcxdu3xr0JQyMWzCxHdauFCW7OnkU6Gdyphp0iNZ6K0LVD2j38S
eUyDA0ImFOcqS/xQxoHHEIUYHp19FOYBnlU2Lye2rWLNJujs8xzEAZu7UDFMSkRycVeI22Fj1D0d
S5t0BG6VonigoORlsmEIELFn4/x2wAqlYB3B1skOsLvB4lRYxPH6gL24fI610xAQFLmVSFZT5/rK
oe4DiYnUmk8mtq4se40Y0SGfkAHEa11QK+/D1PmIuFcsDscdoeY7ESdNyvxy+urY1xj7WA2Y1Q2S
nt+Yz/7fmNwDFYDucq0B+4CwAKzurUn6HhmaS0Ezvst6P6Y/MxuGT0RJlg0Oi2elPp7ZE+qGguO0
2lVxkeA/iX/Yp+CtcrG+sFObmD5JbrCAJo9AIvvaD2RBbgZhkZTchMsRzlYKioNfuneJ5/1Kysda
Zm5GzQT/A2RcmGanT3YuYN/eufGHRgOKxZB5Qb2/x/fWNDBPBBgU8EOoc+jQ7hh4G3l0J5JLUqpc
kMw6m63aEJ5aF29jdreMNIyI0+CM7nn0MUHPuv5qQwCMg9T/MK3634FwrxnkEq57quwvuIl+JLSx
1fwuXBb72UZVgeUGGja5VGeV6oCXAxMu5EjF7tKDE+InfYehajrSD3nxTOUqfvUANB2ORGKDsWtz
Xq9uhQO+/XhIlsguWWUUuUqtDwmm8chipQpOdOL/vNoY3GoviLHHiVnTjrrAWFFMVTtEThk9s59y
iqRWNBhVYBK6y2WcHS0doI/YAal3C5f3JY2l17K13VGz2efRRIL5aW/L4OtqVebwWsQpwzK8LI1i
iRMYDukAdql15AW8vINVLZjNUfUG1EnNWUmoKmVVIFHpYKvlMeZBD9DDQv60Maz40vFP3zsuAs97
HrPi1TVrn636pu72y7htcWursG2/G501W69WWR2Tnxn8jClvNlwMtjtjftBaHVkX5zaHOt87OFkU
SaeVDenTCrUrXF9IP/G8pSkgmSARTMelkcukXYXjS+8rAFoRX9XWYmE9j3SPHIEL+Ydq2G2gophi
Btz0tlB0KHggLLlOlN5IuAdtbSxFHgdDv3afwJh/EXXMwRYbj84GbNmWsloAZXs5MCVmLoBfINB7
F4PnDGzu+mTdLQvymx7ha1CQs026LClUprEtYDYDDAAEsUtEHGjuZS+xz/LPO9slmOXntae/LxJO
AjI3VAVGja7i4+JzDO+9yNASbr+CW/2kbmtn7ITN73PEl5ro8tEASVGKlO1GktM279bWocDjWI4e
2V6iz3sUTYc7RflaA5odzVXx0SpPN3x7ZCuLU+olub8vgGkyB/jMpfGDwLsjMBTMulDGR8eAP6lf
Cd9n3GsSFK0q/HsuInSc1il5wiDma2E0MkvmFGppKlpZu8+4O5KtoiWu2aNTrUZtcZ7S697Yyuh6
tDnrpjUoBiJFBEalPKl/kWy9xQQLa7HjGeSmllZx1cCHPy+n139XMM/IGqJtN/RgncUudiHBynWU
aL6rxEtSzjDcmHhSUG5igAU3XY5VKruvwmAh7v+2bhDipSoZ58l0BLvgwH97ff/LB3Abz/APEjxW
BnDSPQJ3WaC176sSlQ5ebF08j2yoIHJ0ViIpF1uhEPZB49BR5IygBvW5GxT+2i4c9537yLLym1ah
7vAAj8kG7nEMm9bd5ZVTeTerKsj/w1eHCNRuLbYkpTl6EqIZv5jTn2XovZ/BeJA8X+vbiCCLze+z
iBWjc0flMCQe28lgHC7WABDNa4GnjgA9+4W12YfWhuqiDUVdamquInbUTRyJjtjVJvAIhI9uvIa9
h+Z9g8F3P9zdJxvByDXVQo6e9+tqlGif53qgoZtapXi1tmZUr7dLta17ViAu8oasEq8tQBwbEa3S
ouaVF5Otc+kdlVe49LhewrNNGO1lkEMYFAVSQsvaL1gWh3+d3VmiAmcLoQKRF2QBkWLc8JgdYKNv
wwEFgX/997dmtFnkfrbRG1aMBrsTWUW47L1CLE0uKrQ4gpFZTlPGuwHHLwm+VkelG83bvqRTVY3/
9RLVYh4jynX9O9IocjuXIxD97uonh1eCsw0v0UwzzdFnlqOuT02txMWjonj223NXUGr37oZSbUEm
aVNvJSp/9zifToDKx0phubwbr0xsAQuEFfz7mGZhWK1mSSh+RTGxUOXiXxpFZPztSeyAoRif1FRP
1HFISxSJlMBiaZKPzZvHI6ZHEwGrt1QOyXK7J7jSExtJUZtHsVHiRzjLj9+XAj/vuho9+CEU2t91
F2EVTfREtO/1pr7HXJ3jg3QqAsfz1igQ56uWdbnJUKeuKC1ZVtEpzu5Ou1Xj7bONoQKEvHTNSQM/
wlzSfuI8e8zr5xYhQmNb9ehjZss8qe28f7LrMWBAi2jsiHbImVANZ1wzmNOWBDlR9/HFFEabFtNN
4HFi31AHtwfpP1PAULjIKZEePy9djDG+Du3wk7NfKYhISGDm1GQE7L2aGj7fsfDsK3bUrOj2B/de
S7mVHIPgr0ZzskHVBpw/3kNhS/B8UFRBlWVWEjDbh/KmecY31J8+f6D6rROZqgZlUMzourGsNNaX
Pu2KXENAjwrYyvFY63KFLsDcnASVLfkDtyR8XrxEPEo4qV3xrUZWc0Zxq1Xhy37EWZPdZFUM1PVR
sZQ9IpoNgWzDWHw2DWmZ2mjt8pES38uslQhDhQ76R+Mb/dk5g+o+Od0RkCGwgGlHNmbZtmMAbT17
+EtSykKilkWcXaxeyVuWGIWu/GuwCuZzl5LNsbgTKYoPPivwhOXD6w1xf4gh5nIqxlylK2Ydarbs
WjKvo8enxL6jfymcm2CIAUoE3VKVhp3wsXOkq41VQocv/aRT+ANxE8kw4xbXPuEMvduNB5d5IcUh
dpmz1up5qImYE1DC8a84qpgvI+dZ658zKSPxELeQ/95HEX8YWtS4crQ0bbFntUN87wEj+wOqJtgV
zEavbbM1GLLDQJn8UDy6Ka77MfwcwqoL5HiL3qj36wyhbjiVedg8BhqEG20fm1X2bZ6lncdpjCQ1
GGUf1KkXpjL4TkBck6orzxKnNlkE0ljRrJhe/0OzAsLDOkRTTLu15D4VKGezeu9oGwYv6vf8Phtb
sTx4y+HXLmIEHnX4hfCG26tLPqeZCIHhXjk6ARPZuW/kzEWpYXX99b1XLTGq17XFfM3ayfVX9E6C
VE/vA/nDeLcDgcpExOSxnRYlfK1o6wrHDjmOiRt7VN46fDL8qh67xdVdhwh6tbYB+d+4qFz13u+f
xOdxBz4FMLUx0uWvADUhFa8B75f1XhY/MDHdte2vbDjy+dgIYRiy6Z9gS4QswWyg/JPPQ6WP3VYk
xUBWfv8cZSh5BgI/oGufTSudNlgneP2w5YXqdTtW4v90VznifgqozKHrbL1jiANMShYbeOQvimcR
EcjhjE/z2JJy4BxH0ToJ3+Uwrn8+VVHyBT0R8d0sO8SDZPjsKljHpS7yimMmrmzcOUY0fUkvjIqG
QyRMmooKGlAVc48/2hO+30WfznY1T33s4G6ZPlKlc1ZaTN5XagoWmEedx9PROGBLoSY2tZuhWdeR
BYBcpVP1yTTLzG9jlmOj1ktwpOOkboCTYdvPZP6iNCadxr/rpUhqtRgOB6ksyhGPEcF7zewQVvW2
d+8dhBfEQchU3QP9LrkWAIerSC5Vart11APklKcIOX7agxB3NGpd8WOgobztZAFadPlHDGJJTv8m
m00q0Bx9F8FZKdvycPmGWBFKjZQiHhwWgJFG+w+JZsfyt4KyM9Ln4rrMpEpH4eXqkYf3ZyNhGxqZ
2Xz0s8TFq/Gj/h6oLQJoX5ZJmKn/T0oB2EEP6+hzdMEBUlw3nBBmpleU/uzsQtslhEzOUQgYTA+q
9SGwe/g6SmH9fsLi8ntj7VDn7YEnzz4JNNHaN8l7irUNhEMr4RwFemIpy22B4MNe6xq38C6pYx2L
pFswjJ0sySMAYJ5RhezDjKi5WcKxCtWz+haBVO+8Sln2hDdxKYitcOwY9yxGPb7WYS4vq/2Oqfnm
JkHOtzmaH09Cb8HnoWih/nK/u3jHQUh/TaLhRxyHJDmYcBv764JqxUlGiHqjMFDQBxJoy7oxhVkV
5YW/YtvXQU2iu8yACSQ14faDBbgfammN/02JNsrqCRDDnbfK9Ud8Kd+OR9GRNLi4KXrnQDpFWZGT
kNEH0BMROyb9RkMu1UjP5IQePmbx0yP/zVOa1M5Ep3BzMfh9FazlxarVzo7NVTGvBhEzAInAKE8T
1o9vzNS9ZdG/jWwLiqyqL6afH1CIAsvkrWxm/QH7UTfCEd3vEnyzuekhUsBY0mIn6khHq5jcczjv
7xyzwk8fYJhAErSpOfBI7Or8EUCkjK3MzzJKj48qA4toW4u/RLqsmL4i3pTvV5KLNuAaPwInzgjL
6RemB1/6ev3hVy7jQbO1LRCHWsv0b/yLRHgGUqPQI1ILtQjo9SbFgkJf5BlaqL8TFCY4LJ2pkzn6
uG4+TfsjX6H9X3p9bKAxiWiPBOt/UBES+I6qpCyBGXsf2GazoeFq6PGa9F5gNdrOmPx1NIOV+JPO
ApdG+mfRiulBmUA7xeiG+Lh/TzBBZBEbEVgPtJjdfjLUJYKitXqXfZk2LzI8Hr94646or/CvznPw
I87ri2QXgDWu3KRA4aGkop3W9HUFr15rOTp4TZJReOVCo7nr6MFs87RofJ1yoBc5tYR4aNomRjl1
loxWsiyKWMRhWxRgM0ErykzV29N2Y0iPEKAHZgvAMPaDLks5OJ+iPTblebUNiRWmldFiuy7kzI4v
iKtLx5Xv2xeNjOprNj9Vlz+SsMTypUM/V0YtbklZbSxrCE4APz8f4ST7aNkrwMha9GtYKPslJ5GE
3ocLv3M45WK8oNp/LGic340jRaYQhX7LjOJPYznYg6iMsjHFt8LbOCsAm3KP8HY/7D+envJ++zrd
54QDwSriLlnNkF8JJG+47vUulhp1gJHuMoM5WSdP/KhGRVG9FSo+YYLYPjPw/iVJ/zoNZ5+ulleF
Qt8rgKL+Zxqe9Wliod5WP/QL+CnmYjwzJ03aguGvAeiihwmWERx3yGj5ZTEiSFeV/qL1ZEXLCLQa
CpW60bofPUcpirtFhTg9Kjo5+8widinEhbTYNS40D6Z3RtjMFmyUpWxZKMXjIO4bAL/UYWDXWt+O
q/PEyJvk2NuqSS3GXT6Ipjfw0K5GNrQmk1PsDgTY++yp4lj9M3T/314irpbhy9tPA4QV/TrCs9+W
Ve6qSKvJ71uGmOnY2wOmtGEzQMFb9olgMULyBS/tJe+9qahHCvyYlWgH5iZ5mZW/DJfivz+nk7yr
U3s0qjVdZ92QU/0uiHGVT+3uLVqiH4uma8RUG+/4kmzpkNtY47w7zpqyIRQ08qMVfjsaTL5x2+FO
XeJmvOW8ESxJptLnz1XkHn1tctC00yZY/vsG9OWhxsh7+8H1DlU3QN7Dv0A1aWarzEkTsf2ox6Wj
5qJuVBjOcoYZFgiAa2uWddpWkNfZuTdluO3XELc5ZQ1srbkoc1jKsl/V6zJ9dlB6VemtvZxUkNW1
MUlJKAUlXovnJt/BZbSEPeFPWstOfjY2dzeOBKgZ8RmtqDBbv3EPISwlR/LDZzAW25MRbpkOfurN
aRVaVmXm2262bx2WZTl/X7Pi2n12THnTzUVckiQM+zRpx4bNPKWSfiWv1xwLIu2GVZTd/NlWZ3Qq
f4Ds1AQKy4kCMVQ4VBu2W8T2UU9V7wabWwTY3byLQu/KHBriZ6YDGjuiAjOmbKXDw1LWnDMQtJnz
o4r0jMzbSDs0s2tRC8FHLv5Wn9tKrBF3+fwDcEUmw7uCF2FyshU0NUBlOcUSWUT/m9agh1Neeg51
t6xdj3/9ihSSi7XTt0vGmtiMe1C4LluAUUIizk+dyizT1mJB7pf92k50HsIqxvU3MRYS9h2fUb6/
HbeeffGRIhHjcqBZ3qHTL84pewEe3KAtnoH0wDWs+FDL8/6mbIyc+0LSUtSV3rM9ctoXZkh44J95
QJaML1LhVXNlrVJe9iQk003FQvEAdEy/C9CpHXFtLxMJWFbzATfA8GMGsy4XK3wBE5i29LG8RsH9
0n8rt7dlG7pdY8KYyxo+m4Q+BZRU5IwCjaq5kg+9W8NFtM1TvTVQ1ER9UxmfdONW1dg9HMa6FDD+
EfTS/BGyWFyfy2rD2YVM5ALq7uuhbo3cWBEabmPzzVkgYkt8VQH8I7SV60RMsUWAdY7xzn+84b27
jbFD2RjFLjQPe5vHsLHvFhHQkgBtA+deZsifs8zxDT28WABHLs/f60BjF2W+Kx5MCfHO3/gapkW2
my9IQnJm3h89jpyFrXth14mKmNLDJtsDEdajOJojx0urPONcO0FfGrs4pYVvc9OKY+AOcbkqZtw1
ctS922gpCxKlf2Z/ew8f8kDKkpUMoQxXNJCLtTlALy+Ujd880JF70gaFb5uZ6zTDECtL/Rgd5KMW
nGMlQ9Z+f3pT4Abtdi0jh3M8IB9jdpQi5VmxcNwzT8RxoY8KRjEkmz8uRTj/zuMDEuah93Zk899b
R4FP2/knNFnSGMgT2aFmyGlZSRdqPBdnZHeuOejKVCq7B03Sb2gazsW5Bh1rPtqrPJVrrhc7mBqe
DecgTxnpHG+wBBwQTutYnleDeqfJpKcagVYWgmnIxumiJpcuro/p3G50NtB2gPo0tXVohBcMGOeV
ZgrivojaYpMf5EuCET6TnK0C12iHz7DITMMFdCcqw8NuJTPZXl3K8Z/MUgiLFMhJHD92F3fk2XT1
3vim0IaiRcQ9h07d/2N3eG62130p21+KYqM8zRHm6JY845xz8kw+RV5fI7BLb4w77kN6IP/7uZLk
80sIUpsnlwjEup3Lzc7/VjdgN8WOV7nA53tVY1mUg+CLDshh3s7V4dnD3HHlVqy8lqWTzx9dJvJT
V1nTKQ2tfTCsSPOT2DmhKXpWDutk88pHHVDwXNKB3XgkQSjxpi55HRrks4sWujaxtJYHnhmWjPz5
qrPse6nW7OJwHf0BsZlk/Ynftzzu/sym6TT1zgjURnyS7cCRdCUM6pj+1WKHX3/NZbsgAI0jvAPi
k/j6TrGaPdQm4GEuQXsPE0vhH3cf2eXfs3nwnHcVpoMbIaRElcWGREZ7qSJC4JzJOS1Iz3mRWuNK
rc/wxidVNhlv49T63Bc5nnj+jDUtoAEpgzaWwFGk7ufpKodbHx4eJDKRqlyI/cnjVk0feCaTNS5h
Or0NXydEBksOJ2SBQaV5X8vxNCm+MFMqSpAqrJaAuIfXQQS5yAeqpMIRYa+5AOouGxdlwYDOx5FO
/gzACoergIhFmguo3OpX0KRu0dnpunwd3p/DYsmrKaf218vxu/qbxnSjlapbPfB/xGlothaz7VDm
RAVLlkgh66RT+miPh9zWYkO6NePLxKMgoYaasJoBPti/jEMSwhd4EePmnt5kcXzuWNPWaostSoL6
oBBV5Vco4pgPOmlMk0xuZ+NrQgNpQmutDwq/i/Z1hlGf32XEgG+eVP+V5ldTjnWyLwWzoyFq0Ql/
/Bg4S0LBu9sT/lR84dgP2wm1yiqa16brofV+GxxmmNJjdarPXwbin8c7ex6d/YNyhjwB47GIJKor
7iiIAkFASi4lTIjOwI5NeK0nw3CrLTp2tCMU+XWHywvKjqwKaXnIDqYSLvnH1Z/4lHJaV748Ed0D
ra+Wi7r4eRdp6o1+PV4KAqTm6Cu9UOv9xwhdxpklxILbSNWVVQ0QpioAxXU7rnzD1cUbgB8jQMsm
G7qyosT/VCnTa2mct5vm6XsiFiQRYvy6BWztoja348vWsdOtn8h02NP4QmeSYTVY88V3HiSQ7fGU
98KP3JEThkjLYLUWBqlDf9iiC9gJAn0Q1lktZI93uqdZJ3a+UGrPHtdEvbfqonEt1fpLmRrXVECs
3ofuhG8HiHrAjuaTfvKSy2tOChpdo6qIt9CZ6sLrLW1nZ7U8UrsGxgo6tb4JVZKjGErxz6GtYgvd
8+yYOyFvDJuD/jS7E0kKyr7xEb4DjEjSzAJUI11MgskCE2wAStZ/OAWHLKgG31s1UNnNUGEvDPWk
STG5a7Bh6KpaY1vuVcHIIwNPS3WdU2y464ekeNajpF7XfZx0SVMwDxr2hQSYnLMjsf8ZActbsbfE
7DD44x07jEnFBWItzmNt+dewSwzQDf+MKaypFv8I9fukn4FRng84dKczea1PWiKZ8Tu+IuzQLY8C
A/DaxKjXFjGJIeW/xtjg/Cjy/upLlnXDjRZVMxZspusTLHbLol3vwmfZxUcNJnnEqbU8V2qTapFj
NiDg4lojoPsJr5bY4f8F0oijVFsvRTh9i2j5H8I7JtuNNBgndJGuWneTfwT0B+w/Ry9yNtdqvirq
12K9Vr09odaeV49Yu+okMeorWKDsRZOKg+uWZUOcMmuz+FOdz5xukWUTP7+/F+EBXaPsgHwkT9D0
QE58mppmHOLuqs/dllEpfFMNqdiX8mWOEE2CIsBagPbjPlg5oOp8cB5m4m2hvYTizI5bn5Knw5fy
R9N9hu6Bvqtr1WM+cTKMXxkKPE3Nf/9bUS8Gc3gNyjRHbdvMsgAVtZ4A+i8Sm35LRadaqWqKxUtL
nQxV8QmnZrg75naVrHUu+7NU2CGcwOkUvaH8DoTOkgiPGZKtcpij6c8pgrQADfh+r+lHc5OkoREO
nZ72DDwokd9T2VSFWwGQtGh9g/O8xPoEOrhBHhxxTgYn5VKiqGuKmut+DN93iIt8LiDpHHGaJZNG
woY3aLCC9CatdSMJDU0NExNUB52MSk6TJTiT/oN45gH8jwCarwfnEP/Yzm1wlstaZ1RwzJcST8cm
hO7W618f6EZv5r+9r5QmL8KFeAPLS/uPmpsc7E8ylEqfqsh3Ary4QR+FU7jKDHNRuJu2+eaelBGI
BA+feanRu7ZYE/FKV5YObiazvKcMc09uBU4DxURs9A6pYGVUk0JfmSyu3t7dp26nGCN2aE7tSAgu
5Mny/Oz7dgKd2vqu/ZU7VNGLxrKWLDdiT6GNXxZjR7rhS0p+8rEEIVZMQUJpd7XUavgf3C6V22Hr
1q4A82mXUSBNJwXqDqkxCbfbIXRYxAUse2H186yo1ZCpdfthu1clRSoMo+rWTKmaia1eyUw1m3Ls
BBLxaVIEZD0bj+N9Sh5zxPugTdGpgDYaAlmp9UFIxYD9/51Rq1moweJOWTg97uAa3bFJPCpBDLnx
6h+jffSeQ2ix4z7fjhfnhf1XTeSsHBAilcuCNJQvzEV12CumHm4wtLmkZbQ8mB2skTF4rzBx+Ecu
T7cQ4KRWbnKtOwTR12qrdD7UwWoTRM+O/IS9K6wRcBBd/tpHy49VVNhbwGVP1HQReaTrtkw2vYte
UdvfCUgifvvCbUvJIbzWWSWNmiIpGnFVIachyjBEW9qSJmhTI97++syE4FlnOkpNJEZnvXYYJFmK
w2X0oKMqn7G4MZfMK2oFcuDcJSnZjSuPGuxks6cjciNcTOPdqbjBIgypbiIkdR1LYE7OXSqq9nPQ
6PaFM8kSV2iFE5N7cVRve8etn/4dmaO5KhlQFnURWazYW77ewA8irr2u0i0A6xRv5sVRatUG+ioX
ikw9int2BT8IEN58tRSkno/j96WQN3PiVJKfLkP696V4ZwdQErHpIhoYmpoQ5FJkRTfYNgGsKRpd
WwnvDl7wSwTcaUdYDvTBk2rg5N9602Op05hJqpebuXy/V7+qcuHmqkEKm8JLKF+6ywV9ie6tHikg
rfNs8bFeMhSn03kUSDgJAa0Oro8dtbaGeWZqOxm6+Xo3YVOnDgma+nwPJkxP2maReJvY6PdSGoFE
yuUP4fKmelN5hkzXNaUtL20e9ketG0epk7Z73JpdOTRd7pilQyXkmYtvZ/DT8AI2oq3Uq6TbFwfN
kM1agCd+obia+duQNEQ/WOJ87aWiwVhmq2bsYdv6BlkKzCD0S8CQ3jkmQCJvbF/lV8U6Lno3/pv8
2xdnEVurQynC0wCh4ZoE+pg2JONpu5Fte1JRB+0KhYUnfIkhVjsxg7UOMv4oXZo9zw2QLLoUHFG5
Jpm2N6D/NtxGg9oEZ9iqhJSMs+A1RrQyXbhGpGlO1ENLhcTDnVgKInd0gFnVqUXXy5DjPFMfR4h5
D3yrsUo6aSNmzBACCVxV4WqVcRCJWO502XiMdZTobpGSIumi8glGVH1S+sCDIocw8KBBgYjl4Zsw
n5rVGGICAotVyDSsmuTOD4jtFMOJbDd/nMvJdGCizKigvbl5NSNc2dfytEWAg+WwsGvrCInsrx8R
oxsXdd3VI4yfzwghvQBocivrz3dWBOW6eHcSbEL1uQA1zfMnDzdHmg1N9W5UBJa0cXltHqgd0x9O
JAEnLVuX4LD3qVIe8S2E5CVaBNa+HDZp+VA/7q2nWhHP9vRcMjsYDQpQvG3z1DECe1Z1XdH+UTmC
Gppc4JS24SL6LQ3ftOtRA5TeXtNfp/dGPlU7AgUR02eY+BHkDD9dU7CNn5hH2xQ59P0lEyzYy5OK
mdPHlomJzpee4i8YrtpZQKCSwS33acMuAWejmCKc9ZGN4rQLt3F0qQJVoiokGdvvB30mf2NNneDQ
HnjI66E1jYPhqOUsZVUjpHnmVaXlrj3TeSZvxFYYNJGQmaZysWQA4hYC2Q9ii8MZe8+r/ykEFI4G
zP9BAVKXb19GJsDSbGLqwQWSFrgQWksoO5V263/Ibbau1gwW6eJ0tGIpF7eV9isTskCECxn4U0tA
2jnzR04DswUYOZd5sxLUIB92UbPmsssN2u9z3UpIhN36zJKLjjMBX4XagsYKQEQwAjOIDKCBIls5
T+ZUQTcpGSo9EVYLO7DjlUszkq6azXgfPXze8kT8cO4dLC4yO+AJ6U8mYr4dcvnKh6Z4IyjPivb8
U9fESb1jJL70MM4QqH/Uu3rPy88+roI7615t+EwMzj+Hf9/kJdvufrKEodTZKXSoAAZU0kQqNRTK
wq8xBt3GSimKFd8a8CvlmYYBye2iPQNZKIRpePuFE6R0Sk9gNYOetIJM/ekMYaH30QH2gUINwmvw
ME/52H0/tSn4SfjhdUGXvEkvyoowKKGXp49bAH4J5QtO5nCtwXFdvXDU7hk8fEvpiZrOryL8aLv2
fQ5dScpR5zvqHRn0O9wuq+99rOqzQ4GpbUqmZG53c6EUkB6DXCcddRZAWXp3EytkBDsg42F5csrl
lYX7wqEaivfaUGSr00TVLn16iVeDjFLOUyx8DwaNOLUoFi7E/KFVh8pcmOQKfoUfYBxZf+ahJjh8
x55NKiL3QCar81BcQ1B/eRxE0coNMHlqer0mnEgOAmb9MBHLzPswt68jhmgzFvJUJiodd63FFY2y
DfcUpxe6YPiMvSVYQoFNGFalvuUCVBcnItfTV6zvW5NlpFY=
`pragma protect end_protected
