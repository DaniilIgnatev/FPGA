// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:32 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
b1+lS6JNzGaTsv04p6ann1BcXqxRplrnLxUmXIfFnrpM0feUUYBYIafImzncMC1l
KbLVuYmdbDmOXK8dnCZIEcGPOOttZm8MyauNHeYTyf5f/AnMv2bN3YScoHo1UgEu
lGohJN/xUY9cyv2zWhZThxXc5T7yUqL045NO2DWqeLQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14080)
2gsnFmBI+21Yz5QGv4HamjJ1p8PeAWUfo4BXappwFrziGQf/08mYX5JhazAKcHMZ
n82KMRe2YVLEvUdnogDs/1vxNLVWfbDzIDwLeKgTyyt056HeUvS7eiwe6sXVDnf2
UYSnkb37l1eH1Mnb36fbmpmCtG9d4YS/1SFAH7kr3yzYyMIgjKZ2xOj6JZQ2L6Jy
G/IpaIuQ7D++S/Khxy1zK/DlobOz+u+w+6RBYVAimdp2ajuNXejey+b0ZGRpLnEe
RA5q5m8/1yx7l55iVmGBax2OR57vbBHR3f7LLostWMO4yutxcvpOX0U+1/h8TCwQ
+2h4CFteX55x5R03SmqiuZum2IYhrV7OcxbU8uapjxGyV+DK6D5pBiWmq7UVW8S7
rARGiC2cIkniHOX4ZksR+EUP/y7qK2It/J76gQIjDvDgRGGMDa9tK2Nr6ExNh0OU
Vab1osgvZjJ2xbWQVKUh0T06IIEzpBO0afex5tsEIyN05xlr0hMZeAV3adhdzXlN
4ccVPS1/ifm8GP8t8m3ayQvzBBGdbwV/kpCci4bWRq1G57USZ62YFj4aNKBWVa5A
zt5L7Akc8AZt9DJ9lDvGNClg67X3pMOPRfhdyFuuv92reY/xP2Kv8i3hyaM9csjb
Z/v3XuokH3Q5MFjSNY8EoBhz1MorkRhk9+He9Xbo2qsf0jRyq59rMqvVVCVgTBuf
3OEP9uDnYpxGWTnXYUhPy96t2pdXYkL/J2PKC0uAQEFeZKjI4uQRQko72BzXe36X
9S7ZaVzan8POoDRkB5h33L4RHUsgQCM4gzHCBOa6hj4YKX/WUBxW4uZqbXq1Ff/+
m0S8Il9K5YbV6u2Yr4g5AE8N5W7XwFyyic7P4eAnc1becv4P7GD79kQe/QpxnkZ3
ZccFbzM8gDDsIYAA4wXMZSmglaycrMJ3RNfzVhEoYao6wAqITv4MeZcDmw6l9R8e
5NDVYsk21PD8WaGRp3LY4Djl3YLaUjEGtyOLun4otfD6RjlPMrJkJpjms7XpxFDC
um+0HwuLEtqZ6l4CaHkeEer+XIkP2t/aO2KklyGgd/YJCWzqpz1z/4rLHQEgq+R1
4yul//9Li6Td43ueIjhVEuin3xs5xxTVNzvDx/3KbzyiWjDBS5fWRzsNXtxS18IL
kCHy+b7tlIxUbVizd41gaGK9mG6J8btcBef6toWcz87q8lnMZLO6KIUDyLgDpWFy
6dUa40jpQJ0Slv8y5qKsZu+nM9MvNW9aVp/nT6HyTc7XVYCwm8g6nT63JA2y/ZTk
xLR3+SVwTqEr6376lnVDUbGxHhcAIeQFqjKAiXoDsDxktQ/PiNDH1uHthCrRcD5W
p1f7MSFWElRH6Wecgk+QOF3zhhKUyewCQp5K052UObu74G9mAEuU3UxA54oLyZW2
4PEDrehGRkPUUhMA3u8BCZreW4BRq/CGvN3+Be8xU1yQr9/sXVSZPteWIXjJDeup
Weo3j8DiUDMM5WIyv0VLjFuVl6addFPYNydj7/nYVIt/EHomDUGtaIJ70sD2TdPV
kw9H9xTCJW6C4DgE/FYya24xx+GSxN57EVVPos7vv3v4MlWtXPHouFT3wEmrqIT7
imlzUGbqAjmbQsvy/KOqG1JHWNy4swY7UwrP/Eoli3EP/kRxmbSE1TOwwqlI4hCb
0/ir33gKy3V4qdpu4zaqxWrVqa05UJu3yzBa3NOmU5Dn3qe4c2Soog7etQQAy5xH
DorP8Vv5lgW2O7eZ54qnIMNylpcX0loykNBI3J1hVJVBkD2Xi8Bas5erC16otzlt
IDGRMCL1RPFhCSPrzflLM3oA84ydrfQGKjdMLnoBZuzBisRC0RauaIaG2OjxIrLe
3e3Edol7v+7e4v0ahwb5YkZgnL2ps2YMgxNBnSXS/aqYzF03zT6vt1eEFSn/c5MI
VqF9+HjreXxU4wnYGG+BtP/U2oN3fNvpMuWB/GtlbT6KyzYc6w3jAaCD1zIQyQvH
KIJTPPRsg4b3mFxbCVQF9N3Cl4zdJPCES1x7rkLVBbMfSqA9t3kXD8tVJeHmaFE0
kAKgRRe/kb+q2hGYfsj9KL172WbQDsX/Gj9UKsy4Dr0oTe0YFIMIHfROn3nDmSQt
+NbLUHaZYqtMONGC8Hh29jksr42Sq/jt0JqB/DhXC4T9UBquTEoA1YYsJnY1QJPb
WVh7ByseaYC3hawxuCAD84xV22O2AQ1bAiAhkwcWkBIKKYvoCYPOsT0Etn6wBWSb
P4o870lnLfLHTIv9DwL9K14w0+19Xo65cph8jUqNljUsI0Fh9iaVZkUMJAzmDQHr
qjsabvq3D3b++HM6QmirEY9HPdcfqBsMdQtxbv1Q79kfVd+Z3U8sGrvLa0ByK+Iv
vo/5g4LIe3O2zHsmtCDe9usp7cRbzH9oLrLuIE5XZcb2wrCVSo1v3qO3GDU3NFqH
t7TKMcouRRW9XZ00L5gfomyircQEbwBttUKWUBqUyAtWPrjxNoVJCuDCpm6dSc9g
EGCNFjtnKD5ZxJiHS618wzLs0oT9l2jmgUpNfRrmpcg0mtIYx+mMYX0RevKUhrTv
gCous3Op8z+6QBMYR29opuuXjpnO0emqNFkLRcPDoUnh5BcPISOaiAJenTvV4ayj
IkQ5VE3+Jhj8ScbjlS5w9W56SeOUOZ+DD8tTiaomy+1/6asXU5getSugjvS02ld1
s7FOYolf5w027GnCjg9NlDsq/pCGqvM/Mu9uzags9p7grF2Bo7EI1M5tv0iHG658
eBcOGune2Gc5frIrxT+W2F2J55ukP3Ky743NLGuM0XPRTpd31JV67A98n97+oaGa
VEDXlLzfmBsBRWuwaAmlqY4w1gqwA7pqKO3l+RS6mHSu0iISTW6NQIq0a4PQ8cfz
EAdEao4yEbHhAba2CqE5BbZ1dRhuA5MEJ2RWhQQ2nOivd5EqjZMUm9d50QL2tA59
HPcab9aoSwiZaEK8SAdqfc/reBlwvLRcJ7SrkJxNI9dCWeK1dKNye0nG4b3jQ/Zm
kiaaVl60mMZG0sQOuPkDilAD+pLTRPddT1axkiG7LnvTz6ItEo/92/xlqRkkBsQc
rxRAgY3Nq9rrlOOFXUo/NaP8Q82cmuM8XOeEVOh9AUCblDtpyW3ew+0DJ8QcIpf+
oZmiKFFgRWTYK73dTpWjEl59kWuvttpeuNmNsLRk/dbH1MLBqTXHqusfFE1ctQJJ
g38xDQ5Oztw+EyIz73wNnyKafH4LP9mGPMSlMJ5r8qCIs+1gVjxA3qRRixKaFrLn
7dgpFW9uVmDxls0k6OYyzGbNj25kXHU/aHlG+RfKK/YGNDhE82+76aB6puOy2KBh
6i3d/Mgye4nG/cw92KygHUXOllu5NSjRNMmlcH38zi/h0qCtqBUp/7+vrawJa3mg
ubSxTCif2/tTwPMndLwStBb8Iyc/YFZwwOLA3FQvISSo86JM92clvdm6OlRBKBoH
/phElEDZNd5tO/YtXeklSRxX6JKJtO69aWIpMPuzbQC5c/B6WsSGXH4ShB8dP+4F
s7kmHe4TNyshgI/EepXfmj4mW1Q9TO+b7DDu9p/GFwdX4UPAQaSzMFjljtwy80RT
UoI2vIPF95Gh4WkFJsUjeDkTtBvI5vQaqFqqmxapBIoctDGvkjcCeLNJk7ysnhHs
+UCNRBmyx3c1MAA+sL16iBO7sLYBoDAmrQiVn8ORIbGOpkhZUlyh+SaAI/doXtdH
F4YngiL7UxD7CjmnZPBcUHaXOxfODkNL6tybdYql5cG+iWiICXiHwPJ4M8ulhqwc
vwYm1rPjsjLd5axejHldQ3MyA3Jnv+TT7DHK78v3rgbYamjYlHGCcIlSbGgnLz5M
lsxipjOYmvFUTVVD2ykqEjeY2pbF16ghqTtrYgixJUj5eXenubdsh9L5mmlv8qP8
xv9q0zwictjoBY2hUZKdeGc+BRA6IekdDSYCzkhDu/kbjfRFrXv4jY7fjV6UNRjA
HjuMHJI2ZYbe1YkAZJa1dvaNU06YjMPxrEaC5hdDBS71ehT0bPBu56wSdaXi84Uw
OYWfKUHj0x1PJ+3b//KB2Z0dyy83/dQZ1+uVTb24fqW4E+lpY27pnxzf17a6ktp/
ODABrrR/+sWLCQArspcpbU5Y2Fm7gSODVaP8+kwv23B4XWZqai4qmQwV70nOvmSi
b78iobbmDPAKoTLwZ9CRXiwf/M0WZ5bYxBvm+DhEMamD59HithnAnK1Lg6X3pNmD
SOQqJm7RSSOhcs6lMbZ8mkbqQPz9asLHqm1/jgG+JXznoB9fA42+BwFxstbSu8xz
BODDIht9w8BRz0NevPTtql4+XJExaHx/+ZHFWbq5XYayAeVDgkSpVT5N681aSBq5
qiWscyla/dl9nRF3aGqoCtbUJAutdvS1lI0yihxXJAzXG7YrEqRPIqMbaLT6G9NU
67I18f5+PvGZnfFP7koCsjXk1R7KVpjlO/w86eTrfXa3YgFoAQGCE7gEy0B/EWru
UuI7paaHSKr83GcUFpOBsxRh40p0t72Z3D1Z15zwdNksWDNHKYmzTc9t7a76Kwr/
JpSCu4KHaO3FRnxKu5NkOJVJrGvz3nSh+QyX+KAm9ovdUnh3Z2BOzwm0c+mKC1ws
u2Mr4HgtR2WfW1BOM4KdGJ9vsGypmDJ26JP19DQG3YgGCJc45P9fvTDZiRn8l8WC
SkU0kNWR8u4Oclid7OK7p6JLj+Dwtqh0fge//7B8nl821HylbJQpXkMcPUegWkZ3
9NqvqqMkX6p8RMVg9SRd5NuJ1u8bHaiCkiQ98FkYIORk3tlCotEfESb/ESZZbiZT
Mv7KxZ0/wb2XoA0rV1im50qsNn14fpFKOyvzvLB24tIlkJcIPOCnP5Y5sP7yKxmV
VD6NlPUj7VY2mmJTaJUHjKE7QtAB1xj9G4CvqXhvoZFZPFGObaO897zKw/GFJPHa
iX6mpBWF/E9i6WOIr++xCqMTiDvaKS1dyznrs8E6OFO30TYBWBH+jTlQTF5Nhj7p
kl9qxr5MblyKGbTmWFqv1mfrQv535+ADIcPYakRzVDePHyOsIMcZaq1cjSgX7sAT
pNgSqGPupGHCw03esiZJLzJg10Nkq+3itGZ5K/QYvFIgZ04sreMCaZnqDeIlo3ka
Sq9Zq2sVgMlvDBarDt9aNSPDjRpVeAWLALOyauCHP+zKBuwuWjQR3h3QN+d6MP6M
mxXeiMCguFO1Gl8oIfQfTz9WjL/6W4zpAUOSBkgrd5Z0Etz15H3s5uYHddH/AGo4
LVh/6cyLU1wftSCZlzfMW/MUbAMMcxP5fU+Y7bawyGFxtL7gYhxXY1igpUWAfqdy
E12RJYVZihfrl4EAxiUe1L/pARKpJ/IC7hiNWHeoKZFoZGTctuvlNkT73x691vih
O861C4NFYtaLRqftDCbq6rwycUexzTDQUQHzyxBGLsZgZAyAjhGFVAuxkKso1t5E
P/tpZL51PK/lexyrs66qRBEbS8jmmVmgA2MlWEKHuiE3mTw7zWtbuyUORrsRL/67
iuAtMDHQnKfYCz29GXAplHCvYPE0yMKqamlnJLf4IbQo9xFvjLfGXfoXzojQd37F
aiFl+/Vmce5F6KzlXCFM8P+mG8k0J95msRfRl5u2O3PzeHT7fAPxJNP1pP8s2sU5
XWp+IOlL0WjyBERani/qas3xlMP9CqSawzMM8IrTvGxoPTHbAHW0SHhALgu8iP+c
u0Z5gK9U2cagzIPtPzixNGuEDmi7/iUqWRIlChQ3aF30x5lqoOch34bYnhN0g+gQ
YhZbPWAe43lfvZ+LzojQ7+mU8uWhZP5+k8DOAX9xp+zoWt1eYS8NBTLDNb2Anmo4
uD4VM2JwCFAJPCCIiurwCL15JP+dyofkivh2nhL3KiJ58iLE1YyEPzD/R7DIjClX
7LZDrpAmuBTpGAVptkcb5zTUMH16/2K0WY4WJOMNRtrRzpIHM4bWzu9B5GaItwsF
qKEzusmsMGONgNPx8IOpji+Y1LolhKAsNQ4XqhXmMWbM4pnXqPRRa6/N6ZKYoyGs
dpkbvwY/Jza5//1jmfVETR8Zepr1A84OzoDrJ5Fj5OQ7S7PuFaR6KH9H64/cshQ0
KNaHs8vGVgRv8qC975ly30jv9/jI0Bjhap4B5liCC4vzo8SWpqV92G2FnEBhuWFB
Yo0mSD7H7hmbS/HIEWQsZawxyaZpbJKlUJVaP5V+q9mlDKt62SgdYwB9kqFwspKg
dzsyZagqqb+NoxUDkHw+Z3FqXahPjS4sxNJY+4UPbYtupB3JTvMEppZuRMdtjVWU
/YfzzN+MFlmpb3TjUY1EAfCU36AJJ+Zue2CpwtZHnAaLGjtcwkLxxC5gtAcUEh7M
fm6QCRgO3Inn2RuQPcmZy79FkOX7zMJCNeSdnwOcOWVeGs8Jn+UQ/yTB7Ao5Kz5j
I3Eg3T83HilnIvUXGCisu5Js8ZxvCayJtlfhjUyOFhAZkE6yw3iWtBNkMmDZ71z/
Wfp4IqcWnqy68V/hG/pQtAWxNi7WVrh0oO9Bh9NPIzQzSGZ/kZkWxXesffmg0wEu
n+0WFpfUL9wFrLcf69FG9z5kQ+ONUvirfCpeY/bVrdJj5pZvx6WgNZrFbofj1Heb
JBrXrPgEo1ULzpC+CBjGJGTH2e+G/L2du8DxczaPbsCvUSRjpwXLf/8b3oFyE6Xw
NMn5cSQS2BmaMd73npSkrwMB+Hlu+QgmSMFTDPHt2h3BQ+ih+HNWJ6NqRqGS/ajF
nu+mTgb76HFbxHpY4HjoUsI6H4EUiWI2hSVopLNtA09muqcoGPHwlbIQWIodQc8M
j3fbx2OqkWnIa2fbk6wxC31OOPbWuiPtRRz223aUnHY2pyX17Ir7iouWnOBo/edZ
knH1RVfTUh4SNpCb6YZzcuofzJRBWPlZpNyYJnU47ESIa+ytUwWz8lGHvfl/7gHR
LpBAqoV2VeoEzzkZD/6W7DIupdJJWRsF/MvpaTJHh8cW5+BNDwvs8SnLjsTtVxL8
KVQItBmluCQf+Z63WKx5VlEcF4iPhpPbiU/W/amKXYUL40x4RWjBOdRJcghvQt/I
0kJRpXmMnIo5iYw3m3ICLDvHqaBohkDyP48EgAIRAkICxiymA3ivQhhjqFUqAbSQ
+jFngDBswsDClXoRIGoSL1Zndkfdjy0Z0GQGLaNXmhvZW1cNRG9plIV+fLfsGaiL
/U426IQ9Z0oGrNni4BFEFsJAwDW4Y56Gv0KbRhIcDfPRos4+sLE6ziLWVtXkIpwe
2f6ykdTgUMr0Dpd3xlHEUavg7FhOVHzi/ssUGYTtaj5wgQ4uSh49s+HtNmh44k0E
sI9GX6EIYljoMZRgzQPhg7lACFKQBlmdY0IZ+5jNpFP6uIEouQ8iBn9fr5D5hzVZ
vGo8HKjRb/O8uYcTj0Fh67ZZFmeKFWTz8hyG+SrSyo5jQaJ2s5B1I/QV8cMKJjoe
jO6NjwATBLGeN4Mgg6snNvIBkYll16Txz5u0QqNVoLl9nEl2j4rM9nFR2G2ViCMP
xeb/zuE8cBFgMmZood7FdVZrxhTCt5Qio2nW/oKcqnaMcCQlhhM7ZJAGVOxTM6Ry
vfF3OonUdvO0X7JyjjL+G6aNNGjlF6T2EXYNdkyoW0nk0+wWlc2knwvLz1IqnOm5
uEXmWHUgKQTgJ7xYfDMeV4vwRtL84GV6Yi1Y6+FoJvln2igd8lckrQavRkkfINdE
WI+xr0oXjcNvlsJ0A/LNl6bp7XsPZXKUM5IelZROk2GdGLwHJuq1Cg84xzDqtB0N
i52/twjmuocF6LsXJ+q9oVtrewLfGkNm38lcOc4K63YKzEUIFgBLKZxAPkyynbTv
d3f3iYNiX6vggZ/WkuljL9SKryKqZ1bnYn8h7zNeFk6DWdmkxFqBcFgBxvzWse1T
mUrkdGdrqQjebPxYja6WIOsuSSbB/xgMmfQZi8w8Y/xGDsc03tOBHEUjntNrpTiS
wuHHtPpMYvoZS5RAgOkt7YGvgFfec3wmx7Ou6mJFvGivdmvD1/7tjNZkFi2j+sUj
nTiAyE4p0TYQ1xRqNF9iza8s8Rx6mKUpANhxoVW2vHHxSx48jkeNs3fbIbagEeaM
ydnkvmDed8Nty4gy9j3ybOx24dERlPXzwFyMO88jG//uhM5gNxtVcDFdevtfOB8m
bzPcgr05zxlgN77wmb3zSyaU9J7X9rNtH4k9C/otFDiq2CAKpyWInwYscyss5HNF
NjkBGDnGDXHoTi14IrQQ1TiNLfhxY+rHyESXuIdRySOy5GG28+cOnfQG0J/HZzDH
j21DdYMk/MNniD4e5l/Z3qY/ZKqwQDjtvwNA5PRNwhrUqIDjRo78wcTGq/v1AMN7
iSngy6I1BKHNWkmzrsg2JEXG/rrfDabyJnCxOiVXpmmMhmTrPl+V/+q6XTrPqxVl
0rsHnDkmnxdrf4N0KLBMQVYd3ipBemW68CIVBp5kkmXQloTClwAGNTTinU75B+Ls
vCaCMVl2UThH9JM4CqM3qEdcW/TT+EZsWv8R1zeW75bkVKvtTRuzBD6KFrf1JCSe
SKyVOtp0W54hgf8gDbKvSefV4m+P8s/EIRZFwAmF/1iYvPqkj9TvARw+puO8rVCB
PeEZtZVHyptYDcyqf5xpUOzJFGItIshMHn+LGF7G0rZz/pqEyjuNd8Tj1s/Q1APg
UBQun3mhRoHPpddVEMqjMGmTK25sHyYxdJoMfP54BDvumxmDHcVGvQXix8TjFctD
+cDq54VMcYyBFojPSZ7pnM6/n5WhsFA7lUzhRExyCDcvdCc9ss69LMFhocTdZzbH
44Cq/UVXy4+fpYIzK/3uHIwwitxxWsoZUJim5XcXGXdktIiS8TFOCGx+WPcVwVlC
J9js7EjCP5jLwcZgFRWxvvUd7oTGjQQLHZrpf5m2aGlSkLFxhWDJJQekXlhQksSn
+Up0JZ8/D1bdIl2OKGaP9VuU1k003+1eisYWmyTlq4WiPRZSwVjBvuthCsBXMYBT
CYH0xriR5ic9gPzsxpCQ9SP8jvu2QVIT79XS5xCLVd5ExTyIogGXdS9dDFxf6a1F
V6VibqcNppbRUvlrccVx4FPjslLKtz+iJyKj2uOShAc47zPyacasUs0Dc1+rTaYk
wDYe1+yTuNl9TmxY6LV1Zde30nE0Orcb3ilS7oXFyZYVogjUwQ7NjdWknUYnRCcr
M6c6mK6Z8pfC4KBPft583kASp43ogkyoFT+AR2kTtDXYBXZZ+U6ZCFrq5cJ7hNT0
unSWiijUchjtNo+pVaYdxCbl3dgm9NkQhTMCfQ/9/a1EnNSU2xwqlHIFdwonO4cJ
qVwUo+BtpWRQ3S20Ktc+lFQYW7y/7HfnxLZQX/qCWSyvdzTS904TEnmJUh0JWgF2
tJQKDSLK/FvLVVewG3d2i9hDe7btPuTOuV2D7SwX3yphUnCaswzsP8lVJfNU3VQP
bTRowXxHNS9o/OOvOfq57lPZdlXUMkahvT/EEAWFN72B3BCUBC3wzHfX31iuBBXk
Fo8SwNRp9AFAKKZ8Syyc9XKizi8wUTQTncawol8W2aGVWhx+LHNEXel8OlkYhInx
jjaJpxKmiPCh3azd8xWWd4lCeTmLldqyzjlkvcLljTEXrq1RT4xUHzPHPOT0myTI
738FEuP39hd2QnZ0iwWHw3FGDZG74z6M1UQ0kZwh7K1VANz0+7dxR0ThyCajvhnb
FM9leps13BFV/sF6Q4TTjjYdBu15+XgJ1iQKjhrCQQ178qGRxBsXtHBZW0O/tbbQ
WC8mEOnSIcZR6+d0SKNzQZQDfI8+N0WQ/RrQAGXdBOOC1p0bXcU5MS0OHnVHqh7t
wwytGMuCliZHwn3p9PmaZSOfs56Vb2mxI5bWtuUi3qRbtewyuTi2OoDp3807/mIw
GDGIhpcKkxOwi4nGU/3Ho+/JVY8h7becIBXqnjBvDu6FY7IYSXCTNMcT7xUdgqe9
k/t5Qzftp6XzkKCfDfF9YGlamZrOGUK8Na69BYWaq3TRMy3oKGDdaiMqtBOSlS+x
feqxTO9W9C0a7bXJiJztn1oVz1Qyu1dPB9qpnrkdSgk06zkti+WqWP1eVNqUcVGR
pPM22N6IDOjEfXGdBYj1SJb2eaS+2LPrtfm//BHD6BLm8j/+9JhxBITbwI1D68Kb
wOsJK0NAk6UmOeRRqiPi36eTaLn4q2aUhnE5/GlpKCIQqbyokOQ9O7GZwDTrtVUd
h65b3afEF0yXOV9E7UIayiwMGYcYjHpFWp6ar4FfRu00NRt5oBqPImfU5TlnbtKh
S947SG40sAK5G7Jbw179JNCgNKUTIcFEPbdj6JkxH3PuVi1ly3fuQiq0EaFQqr0r
I13ZIOdwd8DamAHlSKmmBIOiXvc8IC0URnPihSdFEUW8ijFvOVAIQlKl0Sp77e8c
p73nWZf3CcFEggv/LK91u6B2NFjf4VFoYTK4Fc+HMSdmGFkrHZp3HCndfAEfzk5E
E/nK8cAaTOkpxeuyK2ZHik33FK48nSgR5vAt8IWeNdPELBjbyDMGMFPXsxYrofv6
1sNSPgZ27lcjrzxgHt5rkoRy98nhbghh1GWrc2tbBNy4cL+5Mp5YMt12rd5xOMNZ
wBXOQK9gXmIkzGQ/SUZLnVzZDsb/0JDNKCP7hryquPlMbAoJXZbpNeNjbyvRh0kq
+hkdxpshocuLHvdAma/X80r/5vFfatwMemiOK+0pljvYfAmDxVW2cY0Z0L8DPnJQ
Fcurztyp+XNrNgrUvZJk8VZkUryIlK5HiLsdZB0VDTFN5EvJU9gh9dV9xEzXQi9V
Le9lmIRRhiuF1PuUWq1/Dn7GQKYI4N8vSm2W0K6j2vSJSKD4N6cPIzuhZl3muMMX
jGmQcy568E42AiUdnoRgYcXO7O72Vl0at3/+JfyaLtYkQieu06HoCdlAwVqn0j5a
B5D+NE1jNgkolUEWOpUHGM57jMLX4y4+IRpSWyw5+K9hhFi4i9kXFRt+Fk07ed2E
GkrEpLE0dbKNbZRue95enWn7mX8SHPauEEGfjv+4KA60zmjQ4f00lq4U5oWIEcqO
678AvkZ8kwh7HmD7/7oSMdewfRk7K+YxfDidnvUfJgR4NoMsLdVHR8tbwM9PdPY9
qJursRXq1qSFbYwNDRvIfG0tscr8BZrHMqQZg9Lyl5OVN768i3oDDKIcUEiYUqqN
GWrBlFGaBXX/OXZsuvN2k27A250SvRnL9Ml5nEmg4acOOJ7Md//pkhRU6M9GN+pq
T/46dJKfQaBKsITik7rheKrlPSs2FweaeAoPbHipoKCHK31l2M9yCbMOE+Qk2u88
siZbePimkcfEZFmRFfGi0ISqtdMdnqzvjUk0rkyhbmdR7z/4d6seBZpfjFMBErE2
J6tW6Lj/CsJm9Dw5LfOwiksU61RxyUWgvg3D4imVhA3CGPh6jctCyuMQwecG7O1U
swa76WobmYZUTfW7rjVzt4btHKM4MwsKHld8uT68QPlVnErpRkY/3mZ+cZDfeRVZ
DOcfsisnTFHRHPGSxJKyC1rlh/xv05pG6w4kupKWbb1S2viUDB4N3RwMKm5iPHJz
tXi1g7mZTYJ7r0iO6GXJv9nXY031+zeTtUMByyIN+E3YMpXt2melSZBmXc9iu5DS
EYqrtcpOJwbQlNKayP1UC9PS3u+mVzCqIJL5r8jJK3saElAnRQV6DadEp9zXWFhw
yFjbnnQ3e+YPnp1XhvJwv/nFCTBvNAVTtXBMbHR85IBzPNlI1v/FwebnTJOFkXfd
XCn6/9xpajm6DjMJDBWFk1abBBRdeEuRbfxdz1WRWLcRNFgZLL4yc8CFTrzxOKR1
Eg2GPzM3TTEHNiosz1hhWlypcafFazYZfySVogo8QmOBrFgGvJxPKGrPLkKTE88i
w30Ze+wKdiZpd0ezOy0wp5jqpGgD+Hq9LvDyAGfp9gcIcBFUo2m9GJhAnrPjncN6
/nTfZSrCftPWNSGXRLNFo6Hau7EyLiX+H4HEQ071a4VbBnIzdrSHnz0536/snhid
R5SOq2ZMSKpGe4MjJpDo50FJpGXPQQUi4BueB1/NnGeh+8Oe3UNIDZk/ZyH0Wg4m
sxz4DVEjfLAG/DKdYgo+2tsL8Zb6Y/mVoVEDUHuZGEYzlN3xZwZTZRGMhrTeQ9L2
2p05+ecGiKNY9ENpsx97hojf/xDzv1eH7Fwe7IfqWtrSx3rwGxO/+GPC10OdWa+J
uGnTF7Z3QgL66zvFF/teGsGZgRqH2a5rUMY43q9MJiw6aCub4ic++ShJLn9yLF0N
3dxr8Z3xshNWV0TyO6XfUJYRq3AKNCRO8B2VMJ1BIueQ5oh79NJAOyhpSntlL5Dh
qxPvKfkWCy2BXSJxKignOP/hGM+slZkOpJw7vXzVJPb2RYpFTO1EMy4J6FNpl1ij
n1pYzU/hTgo9zQukaP3poVM5k0RS9NuF+K0VMAk1oPaIbvoZjqIFonOd6bUvV5M5
VeXhYU5owJ1C/YNRsEFbjs42sRBi/RreOuX4gZSkMj94AIlBxGZ8MEAzjMUdq3xe
6zF4XfpIDjWIX81AzL7/fw956f7d60z5ir8DTjvR+3P1TPrvbQLLo6b+3CueoYmg
KC5piBgoDfhhIR9mUCZt+lr3/R5yZfag7YYNQHuR5FlHU0PxfRHUIBw6BH/wCMcf
xgcPlRLWFCDXsSpaY3U+7bi0E9cyiz9DSoBaJmeBegZJQQUGbwedJihprxpyrvBI
gj04ntuY09RVicEXnnrxOfPj0XxaTbl+FvIp0ZcMbJoLmB2U+DG5Kie2RdLJIa1+
xbk/5G0n5Z+CTUGn5TOS8BP+EMitqGOZG4ssSkyyLzlxY2lNErFUFraA5iAQxpHh
trXFCRcyLvKI1Djezma0XoE1y6r5QgpltTt9AG4xf3LdOmkpGGPGNMF3LkgeemZx
5aZsz1tz/Ym3Z7pa4oFo9P5HmcnbTIFCUgUQC3ZICmW25TPVcvxzgLKmUZ1rCko7
UgkWzTIxqe1PetYaGAb1amoUg+alIToy6Qu+K0peo8g1k4NYrTFX0QqDURQPVv7d
u6HerfD8IUT7TfgHORRXIbt78zXbfv2nth4Ofe9lF5e0QzL0XZayhaQqXbQF6uKM
pV/Ps4AwvHqVsD0Ge4MnNULZ+iBYZQ0Tse6A4/6CuMyJf2TTVgCNkodlqJpCGZCS
kr2L30bxdD4p9MFOred9G8jib24s37xZSzWEZbxZ3pj6Jzz6DU3cdiR/WfVav/5g
u26ULZkLlxsZlWDmt+aeWo9/Q7eIjxWqmtjTMhwYgRnTX7JRPE4Zp+GhDKO+kI9v
UcadUK7nSLfDDb7Vzkt6BY6AwbTOnD3U909vJsQ6jQfneVL4yg2v2/wSCQTMqhHe
Yl6mQdgE1YA3QYkj6lQU/ylOgF6gw/rlG0mXcfkcsjtThU+8NECH1OCPlLYRbuFm
7xTaVzpB+u5i4VncpQx6DZeJlrDnuSum3Mns8D8zou2TPHUIq4dAjn9oTNs5Pr4i
xlKHOVJD6yQoZe1LR8qPK3ENO/+ngU54/Dp/fJTassKF0vkj9KioFiIfkEQyIJE0
NMfpaAF6zVr29h4GhroP9mLIi4Y+dEB808pKMH0Lpdi8AhhtmAb9QXySh0W/GlJV
A0ovbr9m8icqfx9LmwuvlYclvCOx2hFVEl/7KFj/fFu+QDBIIDQmJapjRmzW0YWY
gZuCbVCLLimFGpGHE5FFnuWn1t72G09Gwh3yfCJEY1t9kXVFNOgsIPtrzpztAJOC
Zj+V9/7tiNQyqCnN0i2om2HtHC9iSSt8SQCMFmxNe5+OqF72+vSaodZmeBSOgbBP
e/OtH9oUDZJ4gm9L/s3sOUtgkV+P/CMh88oye+L3U/3YdY6qxSrR5yKtTP82qsU+
fRI9RJiEDsuqYfxugtPuVN4S+Wn4ZcrUzwCKDjjp+MmVHE7smsSEUT/N9Sxs4Fjm
kbw39yBSw51WfFNTvTggUA4nwnSkmduVhKGLsw6SzkM2CSzatM4DazczaSPNyl5d
tfDRHg/mlBeZ3lYkH4hABwKeOM0PLSOGqqVYKYRNvJwPvCENJa8y1Pm89ONK5mef
AgqUbuUciZJFjDZG6M0AjE2qa2O/RZNwpzQVzxYVsdilYRdVAvfbmucizLt9Q9Fn
pum33fMbwh31MhEhgWM6b7E4OOU+goxXpI/mFKCYVFtQARqwTr+17AmnE6j+ItmU
P6iNLIKA+Ro1dIQISXIn3th0bwzOoGkSnQkAOQx4zm26BIly1s31rtehUoInHbjs
+/rpy2qNi/nWOaZLPO2y2VOpr4U3I824j+xidry+Njf6mirMU1J9NbhufuKyQ09h
p/7BniaCXGTdYXNLSozNswtJ3du/7L7LseWGofZf5s7A58IuJ2K0jzI0s20JiS0M
bgsSqzgKomVAhTbNJJH7g80tN4qlE5nuHTZx1QZY4TaxwlTVCRxxiUTeb2GKMuZt
36x0SCrjbVyFZXkO/66ezrmLqMILWeysG/4Oqkhm69STJQCu+MWemEq2wv3/t6XP
IJ/ScItsK7GFEbcX35V413lkpBZ08tpiSgGt2XevW49iUP1Kk+ZUTQlTvSEcET23
nh9H/oyzUyJqiLi7dR+Ndkj+C1rxb4A+JR2IuWz3UZndjI7LPNNfyiVf9rkcDIyL
RzLVaET2aPiQ7+Rkeaew5GxIBY1jY3rf6jZWfp3754Ps1VD88DTKMlxyoBbSUQtw
PJKSsUnpd+vTjWYo4P2oFzzXmLMyWZn2yvZ7YDBQD06whNUzpLxtxZviREEnrzZe
twRnPQfVhsiV20OUwxCzMDm76FgsnVAl3nr/QbwuEfsCyZ9yM8mK7ZxKI9hhdmD7
28jRFFfwyT4SFnV3ScHB9dan/dNzrxHjiciaEe3pIA44xXqCoURi/gLcT+yGb1Ot
kDg60csdVlhG2ZmJwqbzdr2aw9DTfYjul9eNKDyfJTiyBoOOY5N+eAdQ64JhuffZ
1fSmCspfMooP6kWW3xqEpb3Shm2R5bkyNMAs60StW8NtoG821xvdkPF/7IVEkiC9
+LNXq1J+zDPgZiFR+FevmrY0Ic3qNRq/8bjlvVuWJsfPHepSSvv3+iS6YkuVdG0g
Ey0r31xjpX7wMkJBxvgQrMj1g+ZMaHIYuuHtqNapnzbqNBkZhCnKDkyU7iXyGwsD
Vh/xqWg+E7oJyyQ5nhtLj0nNl3dsp8CQdslq30vw7WGtk3CBuk7KqehUD2RJZuXY
QJOk7K4H4NhScNxEyaTvRkfBfuWfR5C2B74qzWwqebymCT0RYZeAjqpN/J/MasFT
O/Eqs+w652KMuHuUxZV5m1DCUIChO86EcoHmyAOk+h8Hq3/bjGMh9v9V/DN96LTQ
k6ZqgXweBecRoJ93hW/FJbN4PBCvhsId6MJ35rHJWVNJXN87qtBGoz+OXCyaYe52
VZm5dCwwihwaAQOPoesjuALqtAzsexD9GM5zoFvGa7qso5zSDupbF8RPyONvDJq9
iMEDqLsku1ez9hNHa9GdzH2zi6BaLcXAYk/PelABoa32MpcPeMfWIo0yO9ELvGOw
Uuh745KsVVE4S/5MJUvgPrMs6rflS/+Yn8VDdse8PQg9Y//4rYcNg7ME8ord7koZ
x+eJTm0GCnqXx8XWzGSaJkGkKc7V5lB63oCisKMfYaqIDVnvvpNYi4erlYuHbiDv
vuPbieQtS7WOUv+suJ0HzclzyogO1HwNQC2SbTC4SbhCuM90Ur7gQgabkcqaHWoP
QBm3opRxXilNFLwNjv6Q1u8uUzA0FSUyAOCgYnmBSW9SEDjt4BpsFkfJL91IsrIX
/M0koFXjMiVjkJTH8P9v/MEIM3n/CkfMERQP4UfN1SfNP8UEYBs2iJuPVYVy9oIL
MWbf1mX8kIMPO51eZTeMUPuTPjZeTpXmpf3og2+k4nhjLYKy/NsMHASoE8beAV0q
ad3KjMSVEWKwh7YAX4GcpxECyCsQzi4DujdRsSy6c4Wy4ZMpkc6q9Vf5xjRXMOAE
UCZpqIb1OVms15HjXkU5UCyKAyxUhALJ4AVr+ufbmw0sN0lcOraKKmocWjR8FG5q
HpFzSS3+MvFMVJk1yJftQvVLhzAO+uYlSA1pAqWjitQr4yKc8bSLAbpGPiIBYbsk
FyTGLqRwyCXJVLf+ukR2DtwpX/Hro5bnEH11EAWy9i7OHX2Fcvj0CLUn/R2q2BFD
g14wMlZF+8KwTQmHyeQLel6G54FmZzq+gKwx0RS3Z6cwg5DZ+OUzNBKcMT/Ahe7v
an7J0mXL5T3QCOHY4G6CFZ3x3z0/Q6O7hh1IczRtdqE+ycGRpKysXgnxAgaBMYya
MH6XYuTTs1R59KBvmo1wMrpdjCy3SnKglylt96vUaeE/eve4mLKAvxb6HhnSdQT+
/xBqsxbiajV9vMl1Ye10nAL2t4t/H6wlUYWyV6OW5OPl3tN6tIKp3X1rewCo8Yxe
uZQTxqGSCD8TJZjCCnichNruEcq8MbpEr1p564YBGqHYplLvE1Sg4c1qNZcKV6B5
1vSsCq5wtKXlPkJVWbKi6bEDnw077cKGfCu2ziYjlqP11QLEoPAcVvjPB6/JApGL
k+89MzFBtvS0bJ2GhUsSpzNPFRdU9LBCJEZFY5RBZnItV8izMgFMBtiGSRciuuUd
4LCUbt0wnt/UifEd9TSJYPynKm27Wcc4o4jQia3tt6ekXhFTCBIIYk8YlHuhfkk+
vuT8Ob90i9D2CePKCCXeIzHhNb7mmMoURsaOqUU6Vbm78b+lBb5ACQwiwBDqAbsx
GJELfIUAPTw8LzCLK9xQutJ/OLePXkiv2RllVORrVDd2UbaKh+8H9kzk8zbioS2c
QvUlhe7ra+c1iKIOV+j/Vceif9UYrwioj192DAZN50GJfkQ9MsdfIsU9I8HHb07I
/Ma0tmSVkyPZ0RLFmLwrA0DeGNmSb1AzXk4XUHudVvycwEB9K+OQE1jzIK/a/byZ
N9tHKVLgSUPCa8uNKmgVtkjaXgIfH4psAT/t+X5BhAm3kOIq6f/SP2mpSCUHsfSv
hFaUOwXVLgStRb20URlF+9Psu/AxlYd4+/9FHpvG4e3SsY/20jIqOMjjeTcNDocs
Pfq5Vy3nTI0k/VjqEWQDM8hGOZq0ZQqwlxrl9kZPmDVNlnIuQpXiVg7roNg/8OKE
qdAQ4JN50C2op50Mfk2LBEdjZvScYWtsqEu/xCk7bNnsH6QSYJj9FoEJ6DtBD9MQ
5ZtO6EBD+gxpTLJNoa6IIGG0eG1OOXnqyXzdfYbqHvye6TYIWnnC/+oHYjHfgbq7
m8fOSxKpJ6JO3ENUp7ZthtxwA2/Im4YbNmqb+IY9rUqak63ScNoN0HzMhWG+oJqM
s5RjuuQ7b+FYFhMc1+yWySJfe7dv8XltfrrBbFvv5gFZD4gtYVk7HW1eIAkt5zd5
N/mj2aSFZZ2BI9hAM7JDeLe117kghGYlLJfwBcI5iL6x/7eYmOGV6FxDOn88Wuc2
EsJ7eJ+BERp9ZxkzA759jzIuphu13O0TW6IlpkN26TnItuKjroPQxxjGuiaZ2pU9
M48RnwhKH3j+LHDVyGB5xU/cu5BjJTuppMeDrnwjCsf+fDS7HU2Lmmvi1j+LxYeJ
RgEzunQ4UudW7CKpIIF+xZ3lv7T8epIKaWd7wKvfxTeSqXjtZYOv48yhrKU8sVLQ
IiasCzsF0A3VDV461J/LUd+lsP/H4MPQX23d0Ex3D1NpM59dV3UWRHUMZfqqWe0b
Ecq5kBv/tMqtI/o/oq+BtpFHxhL9SWG3rYMVvTsKdLwzDeJ4XEplBKO3Y5EYx+Q5
PBAcEEi7082v8mz81uBwMgOl5mG0ia5UfkB7ba8YK7Iwvjxi79hhEVv8l9/yq5O4
w2QXvPqFQMwsieCQN5v1Kzcm8QvNHgiC5U++h80MVAELUmdrDNEj+FV7hWyJoLN9
Y6oC+/XRhRfb0SkeaAsoppFSj1sHg+e0+seq+tH40pOOq2oMsSD6cKS/C5r3uT5C
fMQOlG8TXRz4SIMv0E7MgLxFUGkCOiWmeHJJ6hvHx3fiMH1Beg3M7DxOpf2ZAFcf
rLPvMsRgKUwgfaaGxOB9QIHmrvesaeyqNj4Q0NfKKxr33B2g3i8FYK9vYXyjmdRQ
rbB18xLtzohF5GH/2ipmGj3CZbX5kcLLF1Jby768ZQ6hIKLWHFzAQu/B59v5w+PP
zPzNk1mTQwAZxvwUCRTgr7ra0jfpp699WAZHlxQfCJUBZTP6BBmSbf++E/sMEIGI
zAU9Jpsc2dpLle0oGxqm+MQHMVphi/iXIWcsH6/QyGY+QArcDppE6g1lGVg/RWMH
L6QpUkfkS2+ey+Js5kL8VMf49Ttvn7RVpOERy6Om86KjOCubOJKl2uacdi9D8b7E
4KS5kYUH55VdDEsEU2/B5ilVEPUeFP5yLH6eKiWg7ERLjFZH5hY05adJBs5cZXvU
+6bm+MyXmGypkAiiMY5+2BSPiuwKqys0RK0+u50/pbiIta3xHU9kxM4V6g7BeyDk
NAGFShgaeKCR0dFSRba5CLXUlCLmJaX/Q0VrLyF3BXN1LvbvVVsFPmaxaHaZzMQK
ghFh0vkpYLe1gcvCymoVEuyglaPrKGvnYCWrNcx2WGHtbEkRzj3PLR3EEXKHboYr
hSfJi9hdiIG2obDrcelQXqbG4yESQtT2YLIMu8scG/6lBPq76v45ETZk7QPVQCgy
pWfwff8GkttPF83qN4wmSE/clrwUhOzlETgwe0ytMYL7sRE9vJvxLoAvl17M+gE0
5ywJWvZwcowhrXBq463aW3G4XY/LUxnuE5bNW9cNXvGJFQqnMBHr3FZq5nDf3Gh9
B3RcvNbpp47lD1zIuUE/Cw==
`pragma protect end_protected
