module dff();



endmodule;