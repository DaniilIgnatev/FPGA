// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
lq6PF0DBOtf7WXppPIRdAwlfhkFv0zt3et+l1SvgmDmb2TAlzzkkzu/sHi+cF5Fdw7bTdhDkC/yo
+W97IOJR8zF7ioFr+fo9BbUh/K7eN9wbDDxHN4yK6OB4VoynMeG6ToUkkl0jRlxT2LJjUyh/1kto
TkL1VxglfgYTvjhs4NTBrF0Vi5pMr4yI2l8NdnV15zt3OJSPdeQzfh2YcgF2334JV7yhlDo6N4AX
Z2gbf/1rEetsamO3dPi6IqQgXz+ipV+Y+7eWBSVu1Yby9IrKOxIGWi7vj7JZZEa73674PBZXXlx+
6BmhL5hjhtgoYdkQtvAtnLs2wvj6SccVIpdcWQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9008)
wlI+a9XFz+qYB6DpW+2tLwoRSC0C4lCMMhAqsl+OJisPxGKy8CImkl/pitHJP7YytnGZvXG3j++a
pGWDuDNtMLycxYj+c8eosjkkjNc/zQGtitjkfqTiLNAM+KfluJJYK+7bMHEZ91IKquLiR88sWAAI
qVXHuoXB+kDoGlvvBdOmZfLKnlyjUNo1WujlurLqKDP1O70UPE7hZ3gF3aAdz3N/dnSwwmdDB6P3
Yg2fy3yUDbJYpqn1RngxySNJW2BPTyzLgOWrtP8r/deUXToqqWyglVzOiCkBnz8XBYqaKPk0REIl
Y0PqxS3xPScZaSg+fxnqaC1V1bu1V09vTJhoJ+QUjWNX59qUovoVB9SeQnRvmB9NFVFHVA84JoZf
LdDNl6NaTYVdmOVm7CXlq7CcBd81E2BOU8FFny3xvN9xZ6re+tp9zZ1Ho9uHy5S/ZSy2jyYzWdjB
y7ueeUkrfvqrWf6YgeeIGDzYjmW08Fv6/Chz39SSbQgAdtOYVvHo9l4FJkR6utV6vwp2e7JzOFFw
r+d3GEUV90ThRkpUyI6+Cl+Qz4GNpvqYatRUMh44RpbA3TUGSXUDvcffRncDiRYBLMJxKgJsMPcv
3szhxd/ZhrftvIHvqer6VtQg1g+sBEpC72cmJVIwy06Y7k4qbrsouEr6PAMA60U4WU9t3AhgVENz
fKMbM2UFZ8IehbAgfF6DKpsi//HBMwdqKUOGyNVyoxdRfPOJQQv8YIzosr0ZW5O/jWR1vu4R96DW
aQ2tuOx7b7ZyQyi5QIxZ+qRGyTUaCwhzIr16ipdCU5jIbOCB58XMZ1rPb3AbAPCeZc9KqbhnjtKt
Mg8x/S9Sirhv0CV9BV4c7gyrUBVSuBb4F7zHE7nEMDSxZBU+799VUCuiElzDqetJbasXu8oCEriT
KFZWFJFlYyqDc7tIBeEOQn4SmrP8wyCfgwxjmTCiJ6eNYIfgjtLHCbubcRrip51u871KF55jUp3b
xH9J4mXYHkrHai7AF8ohAGpXoCKuU2wP7wTdxzGjBUu4rtldW2F2x6Xq2ZN8EMlywWCcUq70E5zi
l/7xNf0hEsUkrJLwC7Ghuf0LqLtnSFmD8p6C81oyTw0MePg0FS49BFRA6KLTn8J5yj0d8qWfTPhK
DCPYtiiHAloG+U5t3whPfF7A9OxTD8pHPT79WRgg1zylLmHPg+kNW3/b5zrofUwT/jgUc3JnxXG8
RC+5/sI3DCMusMNKZTScDEfRhGQSncjmA354i4zXr9Kxo1UeOizt0FsuCWaleF17XDh+rf7Nfd/h
2a0DApjvLXhjPyOPJ3gvGpB50eSkgbktTn43dh2SsERU86EvOJwls1NeO7Epks32upmR3qweYpik
evN6zVJvy8UZ2aVp0GHBvkp44vSKGSFa1c7Djw5mdzQKtjGr5k3gjSBZc27ba1jSLKvyhfhZaSoH
oq7Gv02FjPiktumr81+hFXQNE4cuCMdC68DjAepluKNFcGdW/tLTljKOaeoeWUDwgEVf8/WUYYKg
e5kEKj0nZ7ixt3tYcblzvzD2Dw0YDY/tIYlYr18DDKtMP9ZnUUh800eMc3tP2rji+uYNUd4clkYg
DqBySdNk2TwVwdrI02N2BRQqe7hIa6lpGQfPZGRgoj+tf9Dk7RUWbbVQ854Y9ieCYwFFBMfZDPAx
3364hEVvF0/i+t/ZKcId/ez894NdTRtA1SkzW/OLtHC5ckMfcoyMQmxh6i5HqasouLhiNH6CNrPe
e4uofNnbBqLAeGtxmtLf4igdLG0a0RdIDJupOkg0LE0BjlHAxWMx1sypR/7FkYrZKRcT+xShyOli
2nh4LuWnCt03IQVw00xOkzzKiamuyobvFWMnlDnecQPzJe6QRsv9x467S3zLh3uJwI9ljpWZiUQn
LVcCLNYAFI7iUNbqsIPHmpBtQCPbA7Aw45h/uYtv2qsrK4qS2mvqADtxa82FY6iw7m/8QvtqJEda
pvyg2d79Iv2oCegZYMxDIo5BWHXvPblHkn8FXdRCPVfOSy7bvgs5jw4DmlL3XVdSfURf2lMwnFK6
DRvHNf/AT9I9cC94kPtnP8f24CKmdWGgVit2clRocMHNIqYoBhRiorrscHueSTrDa48I0SHHI1+c
sxroZ96U763fzK3VPnFzkOABVFgBV92uTWVf8m4OnODzJUJ6UwHdUM98Cf7GZlfoHUHv6aPExhXJ
dt+9rowAELBFck6T4F+NxaHjyigHEDsGysz+ikzTwjMSRxAIPGBZ/NLbNduh1cDgFY6HKTMc1cG/
lkbiD4KWcApSym1pCmhQeDfuw4eSOGDCiNwxWSEVvHGdP+XqAi/qiGkRXiN2qT4Vh74Ix8/SWIa0
wo1KLanKnsCHR3JvMOq/+xt29z+xfIzrPvjAc3nTBWIPDY0Qh1SP/Ps0Erh60xGpRNVvH844V3Uq
6CuUQZKWH31Z6wWPBGYMVQG2P9+Vv9JlHfdoO7u3Klc0F1Qo3Amh9/Sm/8STDt47r11ZUXyFd4hn
kLi00F8UVT3gy157B7gPj9jnQf84KFOqMlf3j2xoMWUFhlZx0cBf79nPTS7gSsVPEzoU9oOPShFy
mHogyZXSsk8bSYg0nTR8EH9qiUVd4AXjA5S3psBx+gtk8kDrhDC+U0sqJuEQyRkdZIfgF7NBKzSf
FEgrHbXXE+GMoEl/b3AhmVgrputGld2BPFfjCjhcODIBAi3TQU/2rEQag3VADFMPMWRuqwt/UcpW
2pNRD0lKqwgtW5hyKCgK1UudbVSNcsn83WNoa9LDoboIVZNTPPKBJQ+RkAOlm0I+/59vct4a5Pn+
pQbXhn/hdVqV/whtAetiTGjJQpGhXnqoJjBPaZ8tFLsbrNpG+scDxKXShDrMbCkjmgIlCFi8ICEz
/jfeSYtTb3ZdqtTX11XZ0EdeYg4Q8yuko/MV6A26gsdBVlvN8Y+PycBivyTNgZW35VCdMW1xIyqi
+3B4bAQTf9RwqE/X8XvX6Mjd0mnqpWnH6SzutZgv7aA4/4WxOOwrOJ8mlTpZXfjg9YpkFHbU19W0
iBzo7yPBETs58GNPT+fccLKzWJdGGNuHktt/gKXeBTwJjJFxXxWygGkVPHw7vDep/TWreJCsqRA5
eKZLAGRtS30PasjruVa/oTpQ8sa1Vrcgw/b/bZF/Cg92zSpnbzLJcts9++OaDqSVVpZu/P1CZU0B
YpmiwtHhXcRJ/pY5ITbdZg/bYxa11wKmcu0yC6Hk431tnvuUhfRDBwoS6jO4hhPLB0w4DmMPTAd0
VNuDTiE2BeQw0cjmqULQ4565f79ei83ek4pr5hgG1JmRJbw8T0zmBbjiTlouAQFz2xudY2vFAVa6
YQsg0FfPqPpXI1YEXJ26UmrLCtaGXeQLsJ59fDoAq0rqtE1UryXzYIWS2hhh/jpJ9/jBuXujlVqD
JxgbkBzfZd86OqD1UBXrsSTLKwS7JMaC0dNyu/re5qu0lQJin7F2xr5+pUHniU8AjccI6lvGlwn5
YyVcvAo88gXrfteUF3aW6M7oRflthst1gK9EhCQIm1FlWOBniltgurRolk1GoWfPVHVpu8MbP+mZ
VMtKtJri2sCjbNvreAcQcMsukcztWhoiw6Wl6ithlX2fBmnkTlZL72lBZG6mK+Kwr92JAdSFxsi4
qTFWn9eNaeu6yTuXPNBe3z49ZDOZtgi6P7SMuvzE6cHVH9/aDp0BL6H5i04dsmKwS3zOe/u/LbEQ
pVVgx40wUqgA5SRNXyYDIQE7vL9I5sFw64SqdI0ts8BgaSpmTZJe4xTne/gQW32jqCRlcwMa1BKF
uzytfLnx1lQ6K53DMbvX5tByWyS4bdXJkx7eAbrVelQd3nz/en3NtbOLbOk1TTyf4SvAmppR7f+J
ngyen9clDlhN0WiwpjiIWZFr+N+WSHmdFm2MuSE84wyGwlro31e2r+tcywsMnrI+NcRs5dtHcBRR
mzZquczOKwLsrzaALKn2+IAjivapzXwGvYES3J+lrshp5EO5y+3L4iLi10Y5tu0CwlibgMdgrqAF
owQwO3bwLSu34NKkPjx4JD7P4PMdij57qrx0Owvw44Jv+tzgOpu053thH0qUedNTlnsM47bV/BPX
XmICI5jjWScZdcknvBJe7rvMoBqlibZkOykZ9NfPXWcEgESoL+WC8nWEkqQiYmabk1k6F7QYR9PW
R964jchHgY5WeahzUXkUAW4XbH6d+rclLKk9om6OBZTcv7g3AuxoyRlRsTZcoPY/F5LYNdV6hfiS
6hFN49jyWGOIBidysC5759zcYvrGpRvTuh5nUfGPdGQM4pjphi+rs1MrlD9NvqqQQChZqZyNWf9+
CFayMn/OfCBvGC8FkLbKeGcn46HJwF85Q2iWd8ZoKdFQK/1Ck6CDQWbh2V4Zqlpn16otXsThuIvh
GjCJ7DKYqk1ftQ66EpHGIqkZLxgfufBXDBJkJuxqou6KXekQb0Gs0exZgDE7qSNBBV8+rBtSoObV
DMHVNTskUzXewLjkYuiTFJnyrQQ/3Ic968kyPt2DwSmVLtFIiE7cbJnfKC3S1Flw3KJrs1TDJYUI
hFb9hdg9LbWUEpJHid2uBDfU2pI9l+31mVgqNAQGY/q823fHlBRyIoQ73D6+GvsDumd2GtZf2h+5
lm0np8FRMGHkKuL9p3g7w1y/UYyDBPFPJZtm0yBJXypeHSgdWV7WKrRXF5SzgxFVOmGV1DYDn6Ky
O9krxZ/kwzp6XG/R3I/nL7RwL1MzEQjhLY40lBCUjEoql0tFQx34soI8WRev9Y+Eze5ZEehMHMmt
u63rUN+JR1ZoYuTAR+h47hnhvZFntu/tK/PM5SfpYfrrFyr2dKohyMIB6Cx19RFDGkLAA6QDs0Sr
8hyshcPMT0XHdoQ8fk8k7AiLXpu5o2jPXiogIE06mb0iL418A/NeaLtsaaPPOcVHyUOjp5+5tVoh
nmJeEtwaOgYNr8nNH5ILJE4Utk6uo9Jm0kX7PuCrK0xH3OAHbaqsK0SUYEkk2cjuP/x2H/0HVAJx
o8f7OY+v/Ksy7cen4w6xW+gSf8xdLTNd0h8Bo4sdssFcv1NZr4lueFHRndT5BXq7H/O5Rkdw9oGZ
/hxE2a+jPLDuF1mgupLM7qprtCfAx5yg6FoZUoS5jgZERVoYCPF46Cz0RP178HQvSMTU8LhKaFnV
yAoMwHoiz+3KdX0wEpTOib40ma1BbqpdyP5JQpDjVDtddsye7iFFSVCrdVs4wTI/18AywsWnR2md
tWixvlBwiR00FXXxETwpHiSy69tV7eT/kxXq0prC9bZADorg/JZ8ydDc+Uj6Snu6veUrEq0b0HYs
lG8PgJv177ra/XqFpdPubLTwm3gAul+Yx11+roN+kO/iSSGsxcAyNwxYCdfxRcmMaBsnRnTVW8BM
TLq4kHt44Uze6223x4Hrxk2/SQVFbw/dT6oP0i0byqQqWnLBcU15FolEetKe53jI+M/3bNyy/2Ps
se+Ifl2tZqTGhkK1IXuKB6XxauUnh2J9wf2cyER7wvwG8iK+wA/d0dj7VbXas4bCyMmRlcmwSP/S
XY4BNvwMsBZhyun9+G9BW6b+nftWV9iHqw1txAzvMZfDc9yzqpVZ64lH9SoQXoY9B77ZnGI36Pz5
/LByac6V9uIS0mNzWkgQOPXUa7BSe8A2FVjdcv+KKeampAaT7PvswFoDy8U1qpHJKSuLhl6RMF4f
alD5eyS2Be0NDKsKqJGfn+xYi0lQ1QOrZCvhpcGaFwiNt07adlKiW0wzdYEyVGK26h1ilyKBePUN
s2scKkX/LdUptd0gIyCGBS8CDXaED6N8IcNKtmYNwlIFQa0E1LUnVe9EUlJqrCay9IWB9OuSQji1
KmX5yf5opIzhEybh26n15LbiBELu8HMcKOUgkNFd2LCzXARoOnd62MZu4eMkqzm+jSEnQn5tI1Bk
uUazHrT1+jvfmJwgLN5AYKoMwDT74cHKKLYtT1PHem0QsQkFbRSSscEP0ys50STj3iPimM7LMp8Q
SG6t4vRtENIOrbE55vjOCTLUGKRNPM3TyT5cwt7VX+qW5wqQty6poV9WAivY+a5I35/Dbo5aVqSi
wlGLFZmDQFeiY+drzBGYneciMq4VTW/Pj1l8V0b1ck8YctIuWnV/MTu2dnhhIGKrDqLQzi0hRN4C
emvhov0jUSaDBhXx376K6AxJdlkv1C3/+72mq8d9WrAKxBtyp/mmHsIZJOrV87IQnSULbCcvX59N
Q1m/3vQegOEpsNWONKT1Kw/+xGon+ye6v8nno9wcYl0TeqBZEzvJ7YcAk8YetDUfYWh447Q0WRTI
67Yp39DmbrI0Gx7BLfR5mVO+AV4DJCFXMtKsYaEISC/1Q02ySDd68jj+pHbEPDG9xvE9NfMRVt2C
sJECT0SIrR0+yT0CCPuKsgOAb4OHpz2DUqiUWlmYeQv9lne7MoLRI6zs6BD10aShybBgivzlDga1
k1M2XRVIfBd2RmNBDIc8TuKu2CMmU8vhj2sndQvIAcoRW0CquUH+gymXSCOGRMb+SCO/CrM7YTf4
sAY6xm9SY9iA6iDAGREf/WSiyea6zMYj6F530A+IcERYNvglu82tuXNJ9MpFUmvFD1pLJ2GojV2x
JS/bW2GcogvQkvynXIgR01TIiCMvdMWIGeGwrnmOt499sg9DSvhIzU2CjcaNAUG7ZvI7qdmTQu/L
LB+J5vZQVLCYTcqMy3kbtINoAA7EHI2pNjZdJM9RvtXKKk1R+C83kfqTawTi2aQiCi15sfy+YuUV
bOq/kNquXapBly0W0v5WY2LQUJkwaQLdBQd4C/VTUd5TDyyDmLfxn4jq13j/uJBwmvOiX2RgtEvi
qwYFBfmnf5a/vmzEebEaH1Yf6eATEvXpAV1asrfRFg/cTdymJKR8XTR2GvOFBvkyBBWgJzdnpdMR
K+rgz77w6vGM25ODlWHnjuaHi68pXdneGhTQzy6qfqYu7QXBdOXL0aRwBN1mHjYyt/5Cu9+KpNAo
EXqi1ebMR9zTUd7EvdA2TlMDAIgjNCZSBd2enUbXOO6keciG1PJJUurlqZ2Xwll9ERFSb/vfhx+H
QKbFa97d5GcRC1q0ewemGE3XOcPNR+mVN+OktnF9qoXk/itSPlgfWWQzosrfGsHfbTcxGO5bHzlW
klUJ4Teq4qhBAu3gHMy9Y6g9zVZhEzwnH3Nvh3DM4XxXoRC9yHePJmkgaHiijapTOMl7dU/8hIir
zKv9BgIDi3Ax5dzHblRRw0sSmJoWETeYmVhYyjwESkxniqL3CPneA9iUsYpOZ5rD/2TXfPe6SLCN
N2z4p3C8SyImF07mF889nB3w5m/o+Nf0f5cuDCEU8CqgtS6WYKmqT6m0/uiQ8pV/lttbsjud2DJh
6yaF2p9yEKNyTY+cKDC0IF90LQxW8C2Fj3Gbltq0J8qFtvMpuQ3cdPrDnTk37EL8WapAaCyN0I/Y
3Wm6zRBWBobf/+Dj1ACak0DGho2hSe/P1S6NISKeVuo2wu3Qq7z6GAAxxuY7Et5lfug1n2lHCC0N
ea76dzwVc6SQeSYehOtp9Gwq3b6UUwtHxb0vFt17MegGlyBjeu1FD4rBaOHDUpnMz6Qyw+WJUrVQ
utig8Wh+LyW8MY4Ze3vg3n79URpbbCB2XXuEsWIRm/+GNAGi+vAesUrVlC72FvJRUNw2KjKuZnUb
rUpqB7Yec5maumJ85zEVIEs0dbhnFOs6C5yDEap6JNaD7XI2GMc4W5rQLLqhKll0oUZ3J3XYiTH4
oNxkhCQ2eGl0krP3QJIyGW3jax+Hri9UAULdarGn0pd2SLg94SN0evS/uvmTl4YiNVJq6Q7K7YqH
n7LjbV1qQQayEnkd/nhvxc/nOAP63jhcZgMgfYyPlzsbsExRmjJ0G1j6E3gt+UmdOUPP5BXj7Xxs
9/uq8Z2yZya51fmBzoXFEVeWhf1DfvZGyB/LXKHPHbLL/aO9HFH3qX4lSD7SzvoUeZrdp/dSlnvJ
tfaZMqT1sP8QwXgFMYj8cILE9KNmelYtqCaMVbb8AZbzIZQEyTnlv79VdoK/wtQSu4WgVvhJP6Go
lglmC22YsDeev/wNTohJF4jJpEoeBw8vMpaTyr2fyl853tiEJV7ayxvGAHeO7jKwdE1byzL60RD7
Tg54SuOo1PbJg5vzjq34dZLNjgsDOUxo/B9FM7UrZhuXTF1zrfC/N0oTULx+TakXSNyp8u+Vgw4F
VEumoFJg0ogUrrJF8jCTCmv13R6EEtLGDj+ge1HpYzDrazZSQmvlebd4F3Mo93fX4wzeAPtqoyMr
yHFDd4EqpzwgKl0g4q5ZRA0A9uOe/6AKyKGOhXtSE4pbWBrzKP5/msOPNFPkaZ/Y25nDVYPa2e7d
ULumBNYwLMNUTlgvNpIbSU8np/etLwQjKoYypZt3EIcHLOcyEepO6h8vYCRbJ57A1anxhYNhxl1T
B0DCRvibC3YYXZDNDfyy3gltKXDDP20jHy3nonhRGwHE53INJ9X+9FOMG+/wiAnprVgFY6bIZaSX
eT+GuCHVpYsO7UikEhRW4RIrrC3LXxoOPdWb3iFaq/jE7aS8g0GFcStLyzyfQg8aybW+xwTihb7u
KyycKK6J5OOfha6yuwcCfHbXJ/Qdlg8z4/du2GKmZrohPxfaIRM2hSJLbX8uvIrgT7+tDIWPWpnL
eRGVyRlYDE2Ga51b+dH/9+Nwev9+AFHT7xEIm/ucdc2AI9M2pcoWCqHGzku+ajWjQ0KSM3YdwSmM
6ZyNs78HtEHpntEEmvamMRKJznLht45Y5hD9VIhkmi232E5pgE9zT7hSUMXEhMwO5LEhIm5N5b2F
b5CweBjv3caWjy1jo8lzigl/ciIKzmGowttHug1vlxWini3P/6XKI7YrYx50V3iszXtVgn5L4d19
wt7E6wsO4h4Zcc3/gaRTZQowP6DhbI9fZ2lCfEhDtj/h1LWx0c7lpRpMvuJ0de6OaefLmR5NfDdW
fxPykrDuh2yMD5M0p3CgEnTE76yNM7Ah8ykX01XJ5eEB79gfuxJrvQ7w+zyIwDNJFxcpXLWbC9fM
C1lwiQ+nc3y+72FAMQd/u4+QwiqLWkaBWDkANsP3liuT3pUReIyqLCzaanaV9MomaXY3HbKtJW7B
jj4zmVULNcgzhQlaI9mchIFyGLpVyI/ZxjvUjqcJfgt6a6H25CpBJFD0dfx8tVdN97oPSewgKx/7
ysZ/V5X4Omls/3tq0A6KyFigNd3eaxrO+1Ogud7uf2ktQBU2XT7UZGoaj105YBTHaRC0ztKRZmWz
2jlnF9qIQ6K2ywVij27iFQtS+yccuZO7NLoFdcL3KAb/ynHIW5fLmfWMUEEzRWcmHfz2GiGF0M5Q
Mf2ZOBfL3yv5EhWkqS56BXJvV1+e5Ok9secupvKNoc9+qtPRA0lMtzxz6sp55K4fpZ2VlKC03sU2
Nszg7OIOWZoGjU3iOCxNoRDLOrJSA5cGPhMdPA7AsxnlGdasoPqb03Dy5D/Wq50zWu2qiCA6iN4v
Uak8XIkukDyDUcov0/42N5IVC9qG5h5YdGI7C9tofnbTEgQ6ENMSztp/gU/DEQLb2x1+Hv8DAh/h
Cy9AelAlSR3rCtCQ6BRIY2nWq2BNEHxKa79bxVT9GJUhdH/KDyoAinZQNtGHLnKMNYaCB4fUTURS
fCnwm2i8ZjaZeWeg+UKC52UPQDiUN9/s+w+YdB8ZUOewS/xre2cShhFXQRyrHGhJ9e1az6al5CyL
c7DP7AKTR3PB/dX3r2qRfilXOjaIJCMFCfpAjRJuuWXY4bXoVf6K2+4HMgLuC/6Ks+DvQq8Y1K76
YyQNWMNs366eXYXbbnXCr4pwuKKGeHAYIZW2nT0LiqhlHkaEbhcR5Hu9ZDMyXuqarZZ/CCe0U52r
8m+gPHFvHe3s0wRfgTXoDFOly0Jt4kgC1bpjVJQvK/K8X++F59RKgAz5+Vb/dqWB3qtFj0NYyHo7
6faY8yQOsx3rIkDB8igw+WglQHZDPLpZKMuOzr72WfcbBmLExefKf1Q9CmFuLEUIgQ+l/rhLoejX
FUcnpf41qwnroq89sL4TPKpoEa9bUmip+XybG2lFaENFWKqfcJsf3rjNg74Gt0Gvbfv8NW+OGXHK
wCoZ7r1B6r+D+thYNq2Qc8TN7gOE/vd2EKCuSDBJQ6tkhlHolRtHRiHeQj1lITx8gzO70h/01qWS
02zBd8LmFt+A/KD3XPAtl3zUrEg1mbOJUHX1Gf4qa/LzNZd5Oyb6WTKGlAqnqXhQTdrDgXFa1wKw
XPDzQzqkJwtHgcdkHsIfDZxJOmXhHgerSrL0xDGZNiKydK/UHuz1osXrIX6GNqHEORs8x9aczgpx
qg8kmaVHtwLJ06XlwGQ9HV6hAmQJvmZbNumCedV/K86rlbJf0U5NveHY2iYmZ1kmhJSIEvuR42zv
omyEdRX2I1vC+jL7JBxNbwAp5QXA9I/7hlnWZBMJCrkFjBojwbnAw/++f48eZnu8xZ/cyNPjdHQ4
R3tgZ0ilFZaQQ6SBZQbCS9+iv6KYubZt+GYRDizWyjbbghhc+TJUa1SXRZJieYnykPL5e3vlO2Ij
7U4QfEssDUTt4ShPXBBZ52Q83FeMXGiTVce+Dr5XkhRuuxIJOHjwCiauOqFNZTk+kV+SdBjq6U1D
ix1rAShhLN5ldmfQGU0T4kEPqxrhAK2yl8fDfrAeAsTK/kke10Y7c6P9jRaqDrjMqaaGUz/IL5FX
AqipQvitotUuNdry/XpeAVfZiBxjdoM94cB4Na5Yy6c08Pwq1qNEtkRoxa87zbUeVC9ZzqC6rpWm
RUVFqCdq4s9vxib+IXI+q5vtHuTbqxxBWA1GDLTVBmUwoBLvxxcCIsNvqGtjn2YqyfP67jvkKRJ1
5jaqS5SMm81EQ67CaHmhk4z0E+kDaGBx2STP+4HmGxkQqsLuJl4az/I+khpwr6pbD9eNRSDU9Jzz
5d9AZMci1aVXx5xRhJaNcAyBp5B6zF1lHc+N5rLC11Tae9MzV0kNxZ4SikI3uJdO5b4Oiy4WjqtT
GRislZ5rasfd3uI22V6DUCDAm9CkRT9r0sjoeCKgLwNOCTCVuqvw57ywv4EFpOzKeYE3yzMGD6Uu
fMe8PY0krgUxHyFQBBw7mTzrJZUO10JA5hEsdNhHim6q877S6/BXHfX45FaJPRSil75N31iEJnZx
WJJb+o8WpPn+A+2ie4r2zMZHut7v+SxvBIn8D2PjVBM/ZEbnEps8N/OF+ASlmLiRWLYVAW9FNbWD
WzWYNtqzu5SCdnhgL0QCDTou2aHe+ig52iqgQJOYp2dPk9aC9wzPN7SRY8r7U6xDeCpLU+yKpXyT
PqwXdrl7qgZ9rVBlIjnvTpUCNDi1/wM3zSuzD1ntZpiM3l+w2ztEiPwNPXII2UP4YDz0leLajzi+
OeNH6iWubPf6WchPzkfzQ7OTIJteJo8OtLkDBq7O1Ihn4tEpd8ytWywnLfVzwYUG9zLikinN4TKj
GjlQF7pS20nV24CfElZtV8tM0kXcZfCVffoKBS0mnTpIZ8/UR0cfQ4mjFuPU1kyrVg290IdJlzhh
IasygmGxdMd9HVgDb+Oq+zhOEgZqDG9dP9rs/0qmPgyK8w2lXTKuQqkxnMrAMtUeFlk/s6mjZMar
ZnWDtthTwAiKB693Dh7CFbaZPZ1k085LgmsOOkyHCwr+IjngJ9RJ1NwMDOhZeHh0pQhzUYUKGgD4
bValte2SdsvAAJnfaifNBLX2T574pqvEm5yM+f3pAVIn5CNCRrvRKgbH3r/J5QEhQp26Kaom6cID
L124J1vt+jUmlmwIgIrSKE0+OZiqadfvXP1AKeHLGAm60PE1quQH9WDWJiiZWne4Q69tIKQQjTQ2
KK7pmz8PKK2ugqiaAXvuIgOpQOrCGFa83WJD+xt8HCEdIt+xiBg9CqxaHEDVfQWrasYWJI867I3V
I8fQxoNYPiDctpnDlc/Xxcoji/kxQo7svet/2u/ivWtrI56RMvDkcn1YUcpBQvmKCqV41rtVuJrL
rlM=
`pragma protect end_protected
