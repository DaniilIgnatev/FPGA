// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:31 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KWlkYyY/yofr8Hew1eIRvl9bVATJaoWfWBL23zjp8BiE8EKkyTjnuvN3F4PRuwsx
hAv0FzOFdJI5bqFFJ+A1n6tgLT6nsNJ7XJok2BoaoZr63bOmCPzRm/lOI63ufxVC
9SC64//MLwiMBWuyOXA9xzW01w1UtXknpRkU0Boo0CY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17360)
GLHuLeR71MpSwTIxAsmbse58f0J1EV2Lp7MQPaOqduGMAvHUjJzCqUn2e1HyYRtR
tSLJPfpAmZGLculUTUEfUPp7C2xyolfAKhkqYcLGq95BrLYDKhejVJyZlgCavn1u
Wt3ePdJc0ZegHyGKJVnfxLJZDA9HPyJGL4hIVSDnd8M2knCddR0iJLXYmaxW51Ua
nvzaDQNoxS8S+VEEp3AgFIkMEviPokzhMTSV7mx7YJbtGisU4teamfHSsyZdl4CC
AchgVpMg8/OSujGX0525FCiuPp24ml/mKXNB3Ww2MxM5gHcrCEcn1o7mEYDkygEN
5cR4v4/F9wE0nCRPztjuxwX6mY7e8dtTviQtgN47bl0LmiIBBSZmB1VpWYuE7rCA
kC/5MsuVS3V8mPugJZ3S+iHSM3We8RTocvbwazylGoovBc3yCvUM0vI/Zlp1hU72
NJErFGukFQAoVmIZRB9hHsoMNnZgcgLojTWc4TltKR3NC7VPGYz/Vuuyh4TL50O4
JE/ZJ5xqkFsWyWEqRpUayKMk66KHg7MNJdtONLyu1RY8CyoDeAlfGwbzWiQ6UyIU
fJTk8066hzRX4IR8ga0CPgGd3vFR5lVp6n0obENQ3h1wb31ozFpvj4Wvh9N/uyGh
rasJzF/j/Fp6XmH/zqQeNDxh00CscsPhSs/vy28Z6N2hoYhogj425cuiMLukxg5y
m3POukYBoH3yOVDVbPOwpQMK6xsYzKxEo5lXYGVOn4MaHmamjMhSamwB4mPQtN9u
x9peLaw12dRlhmyqZRfVHPMlkL+iBAGt8aoNzymaSeGLYd9k1XsDRiA/OTi0yTFG
54urY+HXhnX26TWOmfw+PfQ06tB8A0ot3PBZcz987uapyZBGUqR0lPSn5fEp4px9
zZVKWQtMqLWq8WyinnVEZGs8qALcbLJhz3zhUqFj0f9D6Brfuifz3KvZEOUFZ2NI
t4d72RGWVdCXnTbERr04oArvR759RynQjCuJNkUM1RJg9nAf6q6ML+sLjwpcpa9W
VaGLNqfN8RlJKTkwSqVkyykGyNiz60Yl7fm8G+5O70Ck/dj0QsN0UNPcpZU3C6Qt
xwUYXXqQT0phhQLsoCPFPFtpz81vuk5Uxebtbzeoma6uWllMXXfrxJov1AuIw8YF
M9YSC7mmKnXNP9OL1FNU1+xnGPyBzt2mzD4LXAef7iuCZoaByiDcbu/nMim2tsu9
rNy9zHJ2FTUB9S8rV06qPSkDv6GkoZIq6zp6zkBywFA1KXVIlYzW2QtLRODV+m6e
59ufOFtcLnUOWLZXQfaYHWKkrob/zjsV9m7YqgHVOS9r6tvYSsJ569i5haJx9Fy6
9mWZYKjGDZrZJ+ZUS9ncb/0KWF/eenl8AGsTYFSUOJ+TOG5dDgiW++iRQKXxfM3i
Ew3ZyoiDejqD0VhOJKnvIzB5dUyYn/yh8WYGTDjH6G1KvjDy/JbTQYkhDY/rIMzJ
dqisLgHX6HFfZdkCYCa22gUnH+w/MITS9bCadDeJM5GD4W/8moWR+oxFo9itKG9l
cznHT/XTrTr8oeXpQZYveSfloI61zeJgCSuToO4fCrtFlcjtnpphI5O2XsBDroHT
2bPAAYUjPoxfVAWn56C6n1VFzccLEcSSQQ9QrTSMm5700YE0UECC6se8zsnkUUAI
0I7n1Ql5NJUGmzSH6ubi9XTm42Ns9LMEHnOtxKi6q6tCzEHoTndvEUp9QaoYKSDI
CS6ke713pG483SLXrzp5UN/rkGnSsuUCO0/xsfbXRxcwSwGrTmKC0xVKmimYc7pf
kg5i39kJT57ZEXa0oHimboRDrR/cuw0K27DbefI5gkg8DlQMS1ehgWouMR4Yb7ys
h77bcmbqudQe8eS6Qv6EtwVZ1MGU+exqtmrB8yjqtqSCMpYFc7d2BvwbJRmOSipR
QmNIG22jP4mve/wCbFvydlDD0Zvev1IjOLbaDOjlTEy44iPTnmmXtjaXuzp3QUUj
VXhUm9y0/hbZ6uOzaLWESv0V2xi/jlWXWqE6uvwyNSdSMo3RgzzzBK+UTSV7C2nb
PZaULRwEqDCzg3fkjffj7/roPABIo15X5kY1ErEtTte5IrNEtbppFCHBcBycMMpW
6affvUiNAzSjOZYafQPXFM9UJmvEyAa7og1rY/TXqr1Jp2IWl8SM+qSoWVPEHTDp
ZxWoypzgH4Ew7jjVJzWBFoF5SMFmI6iIVPvx5yDpttr0iE/846M1BMyRH3/Yumt9
qlHVwj1+EzUuQRoI8x4ZEVOImOYdIHxjLFzPtxKZ+bEQ5qTdjFb9nWHuakZFkCBv
GL2WMjvXzh1z1KO8Q0r7APEgG2RqqJ+x+d+teirDArcpj1qnoyM/wROUaCRikqFk
2pSV1RDF3FAbPZxULsxvHam/6ViB3rlCf3ZMDzrXgVEH1QRenV0mkv9pYKMr5ZE3
bZsJrTOZoxN8Ts7L8KpNvy8x0yjQWdlVXBskrIRfzspHW122OmKx93q0feufav22
8XBc8ULZz9g+R9HgUv+lsZbX902TkJG6hsR3HEhBKAXCE02OUyRzgB9hBMrptdBe
4DJA/EKUHEQg3OwfmlFmatwSETiS7d+EYM2PZlvQOZiLnc26BjSU88Uz3zdvG+1b
YgtS644fZ7H3uCuoXTWxISSNjbJRb63B1CjgGr+3megAIxuzFYFryfuzIOuMP9T2
xKEDPh8bw/jY0Nmb2JQ6BrMGjYvyyJCKSVvFo2eHLQ2etLvPUDr4TRTKFkLh76iY
EapGaNox4Ydtl6s7jwmRZeJVcLhPcWqFeXOILiDdNR9xZIyd5W2LmiNSMXupQ2mX
EZWFz2VrFIKv315tpLjPr/sUIP9EreS0KlfApMXRyPPRGwnB/wF5wYRGUiiPN1DW
8G7g91qZKGp0KTNI4ZBSQbfN3iIkxgbF0a/k+pwvyLDgtJpDC3y440XgR5tCymxe
yLdxknKEC7rPV1MsoZgd6EiavS/2LS6I81eZks8+JPfeBNcgAQjeReSUe2baiTsQ
ZNFXVycCaoChjHlDlrRah2r2W3LUWSt4nC4ETccz9iLJ1s3idydy1zQ8LDE5xKfD
+S8ajq0tXXKSo5KUhwbAzMC00XMx1HAxfou3oQFhkWKulh0AEATzS14V0DNmLoKI
x5AIjXJE0oDp7yYjuDuw7SjKNLFL3mNPn65FuDkpgCMGqALwvNOmr5enKbMxmHBw
BsYxJjw7OolIuHKFS0A/05rc2oLitH3AK1vocZJZc1mKyGTej8ak7Lo5YIKNHeEX
pI3+NYi6NzjrXIiwn8yO9tuci2ZA5VFSus0WmnQ3X7FTtZ8g2SIoqTPM//A+oCPr
NZnisQpjFXUg0xo/HlR5q8wfzKLnC+qJUStCfUJsRLg/JL2+BkCV5JLveakVmuNQ
T0D/ZiIJRNXw9yxvKcF+oWz+RaeI0yfuGpqWNWiHPRFBcbv7L1mH9oD8HRRWTifl
yZ+/YKjcvSnZPrNbuM4HDYN8MjZ+F4thmH7nQiFICZAHCO/jNfVm8BdUsAJogp4k
frkuaTxM+ZvL2Wsabt8ZeNjWDL1JXHhNZvRRGc9srBke3kfNzW25AxL8rDqAnZEx
FTFiAgJTAPfPYR2UixCkgSxYOqFe19L5/jn9lVEbaQC2gcKEuHeWhiUPqA04nbYb
LQzCIV2MEPjFOn/Me9yDRV82JEqdDRytIuhdveJtf/QItXPzu5hDLie2/EHLcYnM
YKe0GOZ+Q8Iwpbk+QvCHbUqbSYKi/KfF5UBZXreYyYi4GcYVS3CyaL2BS8JjfQND
SxPwJLFS4dOOY8nHSn1nk2Mr3s08dCZsirxPQFO3UNZt0OIPBCPnmXyFuXc9l4Xf
cww/jTxvL7lwLd0q/yrUgH6xsEqQ4ZyaBowmmdB3gPC16zu3L9R1+itp8aTwVSe6
Ks/C8SiXz2XhcnNH5FMmP09v0XJ1K30Y4QHKxz9+xdlaDG5D+VYXOlr84cpUQDGn
RdFc2fzELD89J7b+LH9AnegWFoDukCtnrMWBpwSyoGTvHU3zlV4VgcZh0na+ZJIf
qz7RNxd/mNQB1WhpXXp9Zzeg+G3PMAGSIdMuUj+JXeA8eV9CfoA+OCXZjR6NYKFG
LuPEI9u5PqTXThITX58Kv1+aTXvI1lLDeKrEW3B0J0/b7Ap2dVO4IDVYMaQjH6cQ
O8bMwRdAvcbE2eaKd2D8ctD63gbBJ+UK3xGQ1nDLYrKw6ZSrSwcXdpT6MnPjjidy
t6SjZjGhbI8t86N4YWgoTKFEAa5ObAt7mo418OvVQP4oORE73bo+e/5bODkhERXw
v3/svjq5G3bOupoMFSpKqpvQyhWA8I2RoPU59RAuQXxTjm8QzFB/9eiTruqzpSqT
vu5OQEzqMPgG+cn1KjU0F5S0yrlHZRodizqDJ/mzrI9PYI9iDqoKX99G2ADVqxTX
+RTHDlqWwJyapY+wERbxFApqGqAQpDiiJkZ+PpXUHyO44CMu5WzhZLyKu5jjB2UF
gRHtXxchLSlX1eZSivmocBbKqXwClpYpuND7k2ZnLW95A5IKNJL/0uDsXieYS7x+
9+xboHnSbPta/asBdrKna+sXLyiIzuipmFYHhmwim5Rlg5D0TGgjgsimHfPgrFi2
Ggl8UxX6ldSMCGdcOKOmaGUvPiOzmaLVvHy8ovZ2bULIqJUje/qkT+V6GZ2Flr0A
n9PjbKinoc94+4/NGcOYhk9ZL0rmNFm0l0XAJPYPbz2bwR5tmx2o2Ygsh3S+b9Jv
uilDvu8jPj64mAKdol5eUTtNod3wa+493U/r3ZwwdmJP0YMKh7wUOIaQdPzjI61I
V73d28wAuxCkzm04ObQGtm6GxWBgtsRr4Fd60xW5x/1qU1xMQ3LElwmt6UyM29Bp
zu6rrsKIoikGIULrZuw+bCnlPTARAgnMoGuDTp1B6wgsj72oNld4n39hyVRMU7Yo
dhA4LS2GDbirTIkwUZAHYmRWTbse2DQCg4/6coKp1bHgk6ytoyW4uBIDzCnVV6wQ
MPax/O0iiXkDLdN2bsOddhyBShXaGP53Mm4PpYS4A/t1KjnY7g52/wFcpPdBqLMJ
AusfNB/tlmaR+5cuFyISnKC+04zQ1qHiJIjBwseb085hXsdONn/a11VUeL++SEpB
pjMpgpf/gBZfpFse5LUbjimbxDtkU5ySGZa0Cn0Msy6HYWv9BAeIMp2/WGHclHy1
2aPyeAhN2GjT7J1oU788jL0BFSWMq3xf6rINHj7n15Sq1iDzp0D7WchBx4iQEYZN
iz0mzQo0Lnkp7wucCYjB+I5NlRtNuhX5cvPU6S+Q8ZbzHU87RiYmb07SB6xZmnt9
TQ5jC5ZUFTkjx28Szuh6uSxBlK6miMvNP0PjjEB/tpJAZzLAR+2gW0PAfEAb6YIb
DIyNSh2NZsSOaUzEe34Nf/WmwWoxNBlDEixZbYyehJCx5rV1ti4M3uzOY7E0gOe8
5IzywqiH3cE4TBv0H0kXx9eESKSuUQw6cPabtMcRMWIQ7uWqc3ePwS8Is7SwLCCh
91sq2eUd5wxCm1FpoDm3Fvd1BqCVotUqizVMSgrYdt5j64dfYvzmCg+lvtbNuTNY
OsD4pkQhI9p8f5xj4m+ZxlGFSUeNf0CEMJrufTMA1TS8FIdHdfP3A9nqj4uM/AeH
Lkqqi00N4ldKkhbZ12pTArAS9ZzUI0nnyykdd9NKVZIeQZfk8UX/KY939YP+uhGb
k3qHl3Q7soC71Msa9CkkXiVkvLpY/awdamngoSURStZ4JUdh2v7nSMr22G2kaj4K
RBHgoGNNN3gCTC0NLwzRkaVZpgVYBIDCNETxTgYc1IWU3UcvHwqZrDqdP1YBiWnQ
qQP2g7zwHSfmWPF8uEWX1IqDyy/edaVCYwuR9BqoragQkI1eKe/X3l5G4mCYrS/z
5AzruMd2Y24AzG1efTA0gX7ffTIhG9NY6lckjxLYhL6+tE4oXJZgg6ZV/wLa3KcV
0amEYVaC0QjF+xiJrtn+W4alyx72rkeB55q1yGRA1DFfCqzUALfEu1SxSzyS5Vn7
aPvqKTc9MbafJ32rMQxGys3nh5RVawL4IZFf1VBPl/PHK9ddAkK+pTdNPEjJ/lKH
iContfIDDia7aARz0zQ8gnA7pjcI0yemdGjL0rvzv42khpHs1Q+/jHN8cgiK3ugv
/M5ZsieiDic+/kOmlUjAHG2weJjhtvMPM3b2BWpNZ1eUI7o8WpM/c7QaksU3hfrw
fPBMRyYsIlO10xr1x06q3kc8cRX6wXB8PfRXDWrwx11sO+AqGmOOmonYiGg9wFDn
PtvFDYepvRCQ3wAMZ6e+UC6MoNGyQz58zmFEtmwXwsyB08nnPtf1CFaaxyoQSqWt
FJGAYd16yf74vfRhh3MJufmgPQRTu4wAkQHMG1wfUTji5Rxpt3bVn/xPES0GN9V/
SuTrNRlt4Pt1tZz1+NHe5wrcfidcUph2mguaa2iFmm7Bq9OKQVC1z5dL+wBAv8Qk
1kJy/BQQEODais0ComW4ndZp+0JN9PZ30UUNDw3nSAx66Sh8BJNH6RC3tLlXD+Y+
DcCziQZWRB3s7hDp5Bu2KYHgAGiNe+ahSOqag3HLb5DdNSuweClUIFNFXSV+z5JH
CtdrIkB541KkeARKjf60x4mwbGiIKrZPKy9KcmMvxz4gp0ewy1OytOW4kP/4WEQb
qSrfTPe6anyIc189ylDQMMuFWIfkgQWX+CLJ1QYDfshrPyHr+RVIbRRIEPrj1GYp
mOIOOAzQgE9McOBFlmP+OIK5GdKDQB2fK1liSmfhZRKiPRkd3M2TVSilGT7uyEfG
0iIV6yVWStKvjgt55e+HvvL2t6voAuqzxIGizerTpOk07u6dVsKb3GT3ear/Yg95
LXIg8crUUHskeVhsnbTwm3X/4Y0YAXJ9qCom/BcAt+WVNY8u6x8RvXHEWtS+PC0d
meMxDXsfqI1nWMYtj7cWMAu1v/Cpoau+lM9W5bk/s11WZGBHxISjBF3IBMP4DD/Z
AjCkE0l372OlTcFbn4zMdu+/EHhVCx/kEnHTDcEzRscSCxk7W3DR23ZkatrZ4+4N
J1mmWgqSDBHXmH8f18SUpHQ15S32iVcXrCYZf8JpP38XMOZRPoVK02t50tXyP1Bo
2JNZv/LQzjB8PfVcLDnxcsa2DmLnFgliOja2szvt8Df8NYCE5eqFpDkorfgx3bVF
sYkETTVRgdzSv8hXkOcSAHwyPqvc/T3h2cbhPPGtkTeSsgonKHkZxHhuFhUZZhbq
H1N8fE41BgehKtZgIS3UlHyuHkW+g99Z3gs8EoBzYGMFJb71hg1ZL4nFl4k6Y2ll
4bdvPBnkqwlrBm/sCc/9pa3DLvw8vEcP8utN9y+elRJWXoPK2HTGFN/IQwdVrd7N
N++TRL55pWODZBFm39wP2RL1zvqxdPpfApNUSN3HmUMd43ALL4MYA/D+S+m7mPhS
4ePuLtqLdEDVhBsGmleV1/y4VHy+xkw4Az3MXMZukKLcVbBDKux6BngMfBq9FUli
HmllIeAGtCcxC88lDoZzh1m0CBd4S/UMST0Wex/CwzSIq0gUmk3lIBc9KmNi3JGd
LsqO/hPIh+DgaOJoAeEGTF8v41jq48z0pJ7OE9BpjTPaAA3F0qL8vbAoDkqMxq46
101Snvhl0527wd6F0aRZ27Lwc9Td7Mp5LOaOKXmAioL323wu5xfNXa0PzQ1+M+xp
Oy4HlUf7J1uwXrQ6prbiD/oUvvPwYva/3LNYKokB0yhXzHA/LVMttW71FGunnOQ0
flBAyWkp+Ba5Hml0yuvAaHP8s2/5lw6eBqF4R2wOWJYLOWvRAUBL7D0zEXkW/NyU
9SISZio6ApJH8rRDqBLrYXa6EmAmTSNGJC0tgwSqaocMSMjhycNxHrK2tQ0V2B4o
FkNVr+vh/tjvxBAzDxLALVBMauFPRWEfLNM15eVF004J96Z8UCu6WCtsZtifjMxm
iPVngGMDxEOqb72NNQ3XOtQKDtCKSu+A+Jwp6YtBzcgR5lW9p7SXWUCHOS4UG8n/
X4Ubuom9kQLPmpiqoKUt1YIgt3OOFT7xbmsgroY9Qo/IqeTn4aQhIBpFneR8LUCW
sbS/GIO6DO3puFlaYLBtbQGsZLbMdsIzQqZO5Chz4AEm/A+MZIcFj7XDaRj4SOXG
ICUA68Pvl8CyZFYPKOCH0ZwrTc3OqDPVHo2D3YVA7LSvkh2nSUuyNBnsxVKtahHI
7ZSm/HMPlQSjBicJ4NX56AAyAhBgsBXutwtZsFEecGBn9+UGvHjC7tKHD7S6r0ZL
JGQ/o8Au3bLLc1YCmT3QqzKL4CfPrRgw0hQ+6Oe+Ez+hBcJwOkXGA/VnIpSYjCih
N+F0vwoAZWycuUX0clkTXUY/dAF9a1N1c/HamYKkodLNFUuKPrRyPX20vpdRKC2z
Ag4NEJvsOhrT9uAWieyqvjhvqS15dlHGqq40bxWiu6pbZebIWVbj0QokzuySfIjB
4O3YXzYYqaRgEOlY+KRDw/ftfYiIQNv+j1Ip3HOBpPr7kKx7h8C6x61Ty7Ftwe2X
ocS08pgGfYeLe8yEYqtKpJeCJGkCmIIGwSt5m8RYnHm9FB9YXQPyXYAtpvQCFyLN
gEdbiLcQnfDv2F7CKpMdEHH++Vih1CoetcOGnTUDtcYzZ3gGO9Fk2K66syF06EFb
ysdnDWnOzpsN2V8Il7vvQG9YcPrPscUlfMP9XTLEKxVZSi1/+SdanHA+ZqN4BNTf
nhNvlko8xDwdK+jrtFBrJX+q3MdqWHUM5OYlCi/p5ItCj819Q+UxEvcszlpqwWu+
aD4Z0cx7ZZz/Q1zqr4jaTMhiMTw7LyTRBf4SN7vh2+/wIjvvQWnjEEixOMLAdgZ4
a8JbP+4lo6JqZwlsPLfP3zydx9AZgVP6faBho0sCJec+aSsW+i/V0Q7bqBjjRp8B
0F4tK5uOo05uwiBOeEJPK3LsDWh3KC9Ps80EjxLlzq8nnV5FUnJMmzU44FYhMG7Z
YqN2taJuk0Qk6tiXZvmvQzktFZsFqgy6DtaB0Re+V7vx/kL3nEF4lKqsW1Z/28lO
yu/a9pdr2Ir36NHlGdi4G5/2QCBFS1eVgs1zwAG+5uvggYx8qIYhOsqNsg9H2dXf
PUvywUEoaWgYdb/iHS248lS/baqJN2QzN/IPE3Pk7r+9i21ECX/3LDCxXRxDt/Rz
XmHcY1CTKjic9kUe6MmNQTDrCH6C1P+250u0pbi0EFM+ZOjTS49WJaLrb9NC4MJF
cCBAIoCjZuNZ+CpetpeOLUUoN2F0BpBTLZK43Uyh29vwRlxj7xr5zAfogzTWmhct
it1/WPj4R71OcltU28zKfMxkBUySkgb4s3LcntEEkFtz+1pviJdP6b9D1zyzV8F3
qVsniEzKzGvs7qq1voaMThjIjQk7a//UHfAFPqX546TPcdoZ44uJrak95xnVEwQz
5moj+da/lnAA1IqdWHRhwXHFvWCA1XU/COcLxJFrnRLT9fC2VWX4QyVbLK6nCAUn
dRi9udHRCXMwtFVJGL5lK4j7Hf8PmI1GFpYpzf75VjzxgVkvbOebI6Xf/0EMFMnu
UC8C3olZSow2KbpPI3cas9YP8Z5QhVvHbseOHcjhnWm2xsOCG+lU5jLK5t7lTzBn
8KXeQXybcJ52frQXqCzHjCALALFMLQBsjpkl+luhoMPvZa/EYSL/omOXgzy6EruM
fIvO5Bqz3sPYhakppz6wUsQmmLnSW3cKIqbxbOExF2nMG1vuP3cF6h7rtizWW7DI
PLJxlshe3BQqjSRBXuUxZPuKMXYyunNTG/8VildarY5fDQjK0IfQWlOymezVh65U
t8ToJtKsz2dXFER9XTMtShDIw/ebAz4dnMeqtSQvIfxSYiqYmbNCiY2rPi8iuX61
wyK9EjUuHIDmQgMECz/qPJ6vYW9SM9TCH1Sdok41PXACGDtEfxMq8u+s7zlrp1S+
icK1/+8/ibEyEIBAoxHqDb5yX/QqugQoEoS5o33gEuvzobvahACW7KaQTyoB7wl0
zvq8xjj9l0xb+AXbQ2L/AnWA5MS15kiqO0a9Zu9JhQxOjYh1a3AaYg1df7ujXh5e
VktepGFwh65WFIG8TFcRsya7lpnJUc/+pkMsDRSgUZadrezy5ktOID6HPzAm7GFA
K8ek782ZVdS+LwFBiS2s/yXI+ppOod/qHSyJ690ECukPXb4/FPSzPFdbpoo19yw8
2cskwj+nvcPhXhcp3lBx3av49V1vAxCGrgfBSLJn4rOj7qlA10N0vvuEZonLaXz3
GFF/hS3SKlPtHAXUPs4jI1AxgE9WX/yB92hp01Ols54KjzfTOZfyINHh9PxRpqAx
HtSE3bvLgsy0uUi/g51Hzq6Z4ChrQLWuiK5pKbJO1ndSIA2KacHWemMBx4XOi7Cl
k/VyFg7URkaaStC6NjPWqmXnMUQ9x0DiN+jfVEjgiu7CWXOdZve+xFWkbg/yACtY
THHoJeZTAmnHtsCvawgp8Tlw1ruRsCkHWWHcvdvST1DmEZRpM/Pz4Dk7JHBATNbS
Exat4Pjt8vtTVpKgxgAtW2uBQys/qiwOsNlZaPq9mptqHyI8CJG/JqM8BpLEPTVe
s8Zm7APzh9EO+7/k5jhoeDygmstj/LFD3oLrbbLQsuq2s0AdQK6CefGgsnR98o9X
C6qhhk4mkBwFlRGhDi2of0/Zt7uC7pUM6JC6xoDq+ll6Rqhsv1+Mi8OQcihnl6rt
nHAXo3yoA1MyDx9c6P62pYuw0a7luAWFLzm6++YrffmsCjhIvwMJWbgwIZCTFeeM
jt+fSXIk8rYt4g0EiCDbWt/74IC8W8Iwyxt9ivkM4mrxpASCJn8DIWkteRODKMLF
9FyxqBj3HkSfU1TnMPolOv4dlkBYtwWjiLyFgnPCUizoBHG51JiDqXMGjWNa3DJD
eOzV1h6qRuW9ZojdNISrzvImaupnJpp9drpcSiu76Z4GtLYrZcA/9ckwLBKp9ST4
Aze9Hz+i8KhFT+WFkxXaTONlaWLnbgA0/mc0yNyjir8ZZQh4FPeMJgzM+9qLk+mJ
yjjvIGLY17Y22FKOSP+toId21y2lhppq1hE8k+HlkjJ+NMJerBOnkZsowOOIAnSY
4fHFJxFvlYGHaPzPpeYoQZYURpsPcHC1ukLoSlzMAS06WG70RS6srAi1TjnZ1Ilw
K1QrFCaaDXa3AWR6Fec6kBpTGfpY1j3N2r/kt46R0j0RrGenQhWMmlNSlrPaFaS6
2OzQcLPLbCb4L9W62XmMpvXEBVasqFKnYK5VbQ7xsNrJumI1yipDnAJ/32eSW6LI
pm1U7vxPQ/9kL9WvZoTEJ+Qr30wwTP5lgsc7vK7iIMMtTFjFAfwRsZjvAGMy2bur
itr3TXXUkawvu2ikF1pNOJfNrvPN1Z6n0u6ChUbkIv25n44oNtttS8pxwBlqtLnk
mAT/7Dhw9FfPqAx8Cm2Wk8JGSwqCxKASauGEJAy9ytWZkiTYqkCBvb46QFjdPTd1
4TPL/N82G8S345JB9quZVajVc1nV2NMHI7jDNw2gKjM/NSEGmisng0ynrlN91x7z
LrydeuMlsra7HJ4lvDzKnXNNcVrFLpkrMPnsLq8p4v3+8PucCmtj3kGDI7wKMLDu
oVYxpMqfNdY5LxqrD7V2IEwvqMsFtp3FURdT6+oJcdbwlb5ZB1mvMnap6jWmq0VS
y8jH0i+HePOGUGcvLOgG2OaGeG7SHN3AZDcO4gMG0ZeEu97NKY8Vz+iHBM94bNH/
2ozQufR7uXyOcd/J2gFVwsUMEFdH+8Ieazot4uJI5aApG1mhr/FQbx7orL/65Ho1
5GQ51gzyxwD+/NpC6/V11oIEF1No0WiatDjVkYlCUiWzIPomIEZ7lwBpGT+roWsK
HorGeQy5gIMMxDpJ6E8cm7SsnUgHJWBlczMHcuTByCNfg1EKW+7lKCB3rGRqilR7
QsMBLkkxUcjRxA5kZESl3Q5rg1YAy8zLzO4bJ2h2zZh1rGDCqmsvvzaNCficXX/V
Nf7ywAusgm53BleN7h/nIVaYB2ZfoPvLQe9aJa72voQm2VVDHSn7RPMb5OcvTKBK
d2+L0YC8xAS8feJ5o1dNiDiojXo39Y+7CXlavpbxStQt9H6VoTvTyyeFG0EeKn6p
SesrV8B3uq1nzgE6OB8NZ4DiXVmUipu+DCzBDP5dP37y8FV5vLJUixpH/VoSpcic
3T3uqWeqOKf9Jclhr/k6JcXXlWMe+O6E0qh9LB0uiBlqChT3b+x8YIoIRxft7tDt
uFW1S75dCYuuBmHbfPhqmPTY49jTE8fWTbGroi/hqncgqU17s6pPRkeSgeh2TtJR
/EyxRgkRKfyDxAXYpbotF1n1MdCdUowuPKg+6kk6a1M/LF7Ae1JliludEv7s5yLm
UJJLQ3/I49vYheaUvC+q4H+dlJ5TBCNHFU0Q2p+vFFIpekSbQ3tk7ScS9xFKKygW
pJdvOQVNzmr3SBU2wWOT8aeWfNEdBFN4322v2+aZcmQ8d7OQ2l/LCRdZPCVr3Z0f
W9LMEGoPPL03Mh44usw15QRMHrI83txfmc6Bz+xKoxmCjQfLgZ3bR6dtNKfpg2mO
FxWiLlZbLZvfvn4mbPd/EbQYWSbB1N70TKjAxYkF17IZkbHaDCKhXIuFz5vhYMvi
ldcdLzX5xymTBUQMgE07AvTbTg72u0wL3Tzw7eh9wJwvXYF3JOIlatFibY4mreAS
rA5LGuoRi276oQ2CKgTtniEpLyYDjoU1FE405avrvynShTdDXxmntzyYow16IRdl
cvZvTYhYaKVmAvNHzbmYbjjbixG/MX1Qsmw5k+350bQlgmsGudFFM8cqzVX18CtQ
4byUnmawMpLHhJMwM8YBMZEcvjLwgKNwiIVdXrJzODQ5gUPW5Nw5x8PHjkl6cfCs
mLsOpy+JXghOxelVj1zX+Av6ADju/nn6NjUrKDpBvBKKBO7sX4/VsOiQjig3zTnz
Sp/ZZh1omgME/t3qAHoozs70Xb8w5kZ/fMTnvHEYMInf344qJ+3fP37ZfVPplmMB
v5+1Qxuqfz/q2fumXN5W9IHJJX0m5AFNn8glIQzDkes7QUbhbB8vEkqTK8nFsZIh
E0RvbyBOIr6dMJU7F5GQ3keGhB17eVSb8L7dv74+HxiYQMJHioFvG20ag/5btNtm
az/iX75FTiyizbzZvD/37/gBjMaDlyicG+XZpxLgfuBgNHwIF7HmGIU8q5wfxN7e
s/LYchCHtU/eVswN4e7W9VIk+sIxpSGuGy9EY3hvxIJbFYIqm1HFsxX4vcqHhBic
Rstncfrm++opaPRCirl3WThUBmRnZOLV3+WE0zhVqdNtNO9a9QYhCxZeBBTYillP
0/9l2hGuAKhK7fYqLL8NQMM2OW74w1D7AxCHTi5VnsXV3y+rO0wt0vSmBdERFz9G
pzc/Xl9FFZrbxdClnP9aLIpnLcpldu2TqAe95TIptqftuq25RHcZ43IEDAKsmoXu
Avw1vkQuQzF2LQUqS4+NYbjeeasptRqskBvnLPSvKNJNgwTRnR8j5pWR3cYMb63K
gbb8zBywAUzX7y5OMq2soH5Pl5q9TRHg+pm5Mc2owKUf3ia4CzhcRUJs4OVRpxxV
X4cG+AKHtyd/kf0mI09u5z72YWkXctWhJp0JS0uVToTkLaYYZZ56rKxFHkXzGC0M
Pq4Egbb+d5XKxBlz2wLrvTG24F3u7pZlvjw9Lsx2FsLgIf+fQakI7CsZQ4r9OOZK
DxokrwtPjJOWOsT2/kfWluMRehkLAAGrUSiAtxWjTXH3yoIa4nBcHrskqGYW6mIK
OO1LY/MbqW3VvAKrwEqz9UxXK7A/4A+S0HGyVWIDE0SqUUefM4e171AWSJiZbIPl
5vAy/Jz+xUNKD8JJQBK+EvIgZ6SWipXOyWn51O17bTHed8uowX4xR3oa7VfVTYoi
An6Ag7ukINgI/SaMk4oa9hpOqQ2DtAvDvgbhjnolL+AWOfbjsH2ZKqbGGahixJig
j4WQD96ux4ey6OAXRiXj/3wjSW5LZPPoJzl+ZY02p2sjwdrxYdNTTyjlN0kqlNrO
Cc8wAn5b71Qb0ThfZ122zG/+nlaWbHFgsr2UCftCANz3F5znLSfshvzRWQED2DEH
3xk7owzpgFV9W8K/YbdxYpSDt/UNwxQkEiHEQ7/2Ym0h4oh4xhabXzSRs5q3gRF6
y6MdMzfeAG25mJJjVxAl+L5ydAaXoC/3f1y35V9YrSPhcvhv+Gq5ilt9pNHErqTo
A9AboI87rQXbf9Bs6paKMsrleiDH87UioettaiTLIESEHZkQ0coUhqk3TsYwabdg
Y8VO+IrVlrsE36Ji9bYvCdzMDrVbSDoKyO4hnu0FYMxPmCKvYy6cAvmePnT6aZx0
xhmu/WU1ndF6BleexhhGOOYMvDQ7VVYzTR/ZfgP0IQC6rUSo11HQseRJ27HflEef
JQuI/6ar+wVlMSzeM9c7rvuEBwLxovPLPDJ9rLF4pQ4nW84wM3Qdq7DzQZ9Tcp4t
MUZyS6OZUntpRhH1d6KmHjxX/GSw7ZXHgT8VdxJ3PdhIEZ7GghlLKAoqkXobWlUm
7IjNfU4HzhX7Y+UmEg3IqE352nm+HQBkVPotGeHCVGfRCqv9CvMK5SAedjvZcxjJ
uRKtnzqbBR5GuCfAnjoLchMSLqlzDzr2BiiSQ4n3tHbrZIj8DRn4fberccsXiltQ
qJI8lCLCxhGQ0sdCbPD3395DAjK36rEYEOFfmL/OwLzTpDAGb8qP1mQD/G8Ci+q4
LneQfydHsPd/0RSsXD9pdQRXYMQu1Rihx76ixGTFI/1XEF9AAQ+eH+P3Z+OESzp+
rvanpdoFLfJblnqxbWqACEsLNdTDog1FuqvrM0RHbBRnG0jSEY0Y0CtW25/kjvY1
Lvw7xBsjudJv6bYiofdHcaGoNNgl08jUmxrNPf/wGRcThq+BbL+hwJHBs/v+YrOT
PNDR4rYe+9gHkAy4OeuuY6B012fqTKJtywt3UnIdYSmBuhNi3+fFZwBnrhs/s8VW
RggRdpFLZoNL941LOADFqh1pCvVBHDj61khnHyellou+aE5YwQ/VhYwC6HiLxZ8v
yRg1GQoqmf5LkgvNXwqFOaUyB/VJxtlqpxf7FjeTr3rvKOWmfVVyv07RB2Pl1zEB
SbXsQ0emZ0jUAb0iv/ggyeGVNGpkeLinOf6AGaWkoSjiWXn5Vff2KojqFebSSGZn
VXdpCvsHWcaJAiULrrbF3pcVJ2kyY+Um7F3j/RvNx/QS05lQVbjSaHKF9bgcOF7Y
B5aoqwxdPOuGOO/Ong7oAcH5xeOxQVXoF33szQ1ARvoga0Ls9RJgKb8gyANVqxZp
QRVVQxT+MAxBe7UeXqs3zZNyV8w7H73DF3h/rpnXNql06v0ZuOqlUuy4WVa5rjUk
YqP2rnmkygUHMa/IWMj9NGJtc76+nOp3nk4AUCRBoI+t769jIiaCKP1xwFonCq/j
HIm/hqlAuM3y34eLlM81QoVJqMjP40o/H3Zg+GOiezPa80lk4gAQqRNGWV5ualPj
uGtDrH93cYhDg1trvjnfM9soZJQ8eb9c7Iav37hAQu8o3FL2JoPG29P4VwISDIbo
hR7482sOO3Z7Bu2uiSUs+sVaA0SkfFVxyx+ZoCzuBwjLvuFZ631tXUv1hU2RT4Vo
iZqTxXroSZmYL4YCuBMF++Fur7buKRoaIr/FZsCjJwrUNMnYV830UALCDfoL3+gR
XHfdtmdgnEYGdJQueSKtuM0aflSblyJdGDRyJuaazTmX6LSbwquKTn5zQSEoab3T
aPcmzHvtXQCEIG3DJMah7krMs7LRvq0OhDSgQVnVQVHKjvx0kXiGOaK2eS5OWF2i
K71rXP+eo2IfzDJp/gNeqMyb7Q8w9ykY43ZeEqrcON3FxjtFvsPN3jNpy0SCmLFW
8jfjwVblmFrHMJIJ/lI54SGOcHjbqpk5lcxwuDsuXs0R76Lo2Ga8V8X7rIOZDyUF
nFJGl+3sJkdMADymY9aQRUS6WAaq39a++ho6DIcUmExWA3pn/JDK/lrwj37ZzrC9
JNrN1gVHG/l53ZQfCRG8lICA7NgQnEGvDG0dc2bGyiL7/yp+F9ymkAf5vinjgjTw
FtQLFN6pq7iAzvjoX508+TkHDc60y7Bh++oe6lYo65ERJnsvTtgMW/f0BNCpjIn/
tkpdzSzUwiJFuOBVZHitnV6PuCEaN9B7rsjxsv7UrEzfz1pSlW0rNZ9JY4FNqYZS
+PzKpdLG1xbbDJbZxeD2okyExU+y5WbJLv0vKX1yKyFHrYl6n53EZMaWn+Yot5rx
vz/OU9wAdHCYa8/J2I4bR5L/kTssc63EXOepjjXu/4Wfso9DvwjvQ1vGgB81opyD
P0lDiu0/sSnBn1bbFiqkyYoR/YLTQMCUc9SVdmPVKx6fGyjHg1krGfkiACX9wmq0
a6qmJWrr6nkO2pNx5ETNG2miZ4SNcBkgd7W94zFhpct4ioBw7ekJiVDmnCzaVL/d
fsbpVP9rmlgy9mrkcP1ioYx7HTdnEAf/dr5Vf2v1LL9O/1sOMonctrlfmu0XMsQZ
9A+Bjt1O5y7Wm5XHHyBq59OTDwHKJ51Eo+g0TMxhaoQ4Q9Je7CjqXHNe4aqewLPE
LoCI2+dq6fU+zmuHbUkGTGZNRfdk8eF+fVhHZ1rSKW9SAyEfD2RZR3KPURhbCiB5
T/Yqhb8+p8dGHk7Xz+6Vp+/qCT9EQImFvugaB+RiKupFUerIpHNGdxRmTb1RKsV2
gb2e4Ra6g8gamqP6dG4xxb13z/PNsNx2x3RN7OJRIGsSnC9eg1Iv9vGWK+NvMhJc
WTtjC+8SJOXdm49hYEz096oBtPgsq8hIzh3UfpzFCxwHlTWbHZT3NEcCKXzii/l3
3xCEbRRGDkELtKcJN7K3tF3MxBD/Rb6OLwiqD+4rNR7xLCilQpoOPqZtEvfZGaF/
DJxkHqu9KS9Ry62WY0N4x5suz5Y2MG4BVHu6rkqcSiYRD1AZ5A7SW/Vtd3P+tX9f
tv23JTCdxDZuek/boRj3088hNsYzj4O+/nQb9DzWNpYvpcpNgJ8uUUg2iL1hUPSO
kjYVwrqTSDuk/f5viO1Y8oldp62w4+XW6nkd1rhbmmsI87IQNrGbwoq2zLkWWoo3
GyClddPU9CebUnzCZB6SvwReD1frFOJN2sm4+mzn34YpN6mlQtZ05CNqpiEzqs4L
SWkNquXuFFIh5xy7swE/vmZB0SpNKzCCHI3wxq9Rw2+5sAOGS0gaGAsI+4GOYusS
kDFKrbfP7WyDd1Dp/Y+t1r3NQb2hZHWhfqvNtVceUOgWZZTZT0slwsIhHmDclFhR
sc5qXf6PhySbvsGNwMTKt9m4qsEIbvpHLTiVGY7CNtNPK6P3jOF5Ea31EdP4eLTN
N3c+Cifto9yars97Y0bq6G7umL2xolxnSz7OnGRgCaTiV0pLcC5l1d9LZGpq2idw
hM3zjTzAy8yKTCBU8wKWP6kUJRH6qCbA77EwfgzLKRKT52SuUgEMXmVW7AIdggEQ
0s5v3rDBCIKyf8IId82L/SghSY9nuH1lk7sLqALIfhUdjh5eS3EWqFxsjCuCQGkj
sY/E410T0jkqdOrK3z7/SNT+ePR9h51DFRYZQ9kxuMoNtC1Eo1cxCeLnVlXEJYPA
f6Y3RfIbLHvwVAISgTbbHZBCaaj1I3dRPoA3YILDLD6jDAuDVfwOpqbWmiiGd6cS
fJq8RMBhLW2x2rxLgz0cWl+c2pGp1pCMHFamF3NEsE+VgePW28XaH+LlctsFTRxQ
zQzddHUg8n5CvGls0GSGwypy+rgN6gQq9Joi1J1vgW/cVI0bPvzvM0tA+W+yMv9d
BSWWsHLUvJVFij6Zp60Z9iY/a/ZcqB1BVmcjODQj0+c6Y5eAOfl/94BTUc3pXSMY
WscKifNdPbP+ao48eK9A01MXx6sOKnrQm2fCfZaSYFEDcyTTRKYu2dfVsWtu0CQr
sfHYLgm6hyjDqRJr/HOy0ZmvYqRIjG56Z4YdDg9X8L0LEVM7iM8aZP54cwUtbull
kx1ivouZT/1B2a7ZeN6ir7W3exRymaHu9YpUiPWoojfmSaSGIdfXjxdo4MuKZdu4
4S+ZyTIlhYH0RrdKedKUJcUgaaR8nHA8Th1vg2e4SUohIdUGrX1evI/ZOtFFFA7n
RIW+LpIdx3RthdyWkLolOIlfroNG666JcIcNGNnNRdK5evAnAmhy/XH/cUuUnGhz
Ok/7IbGMxxtdQ4lzhHCWgIkutEQNId6MpU4bN7VkcNtrJvXVBptA5CI3SqQZO83e
OIRsxdQDg6dRzBnP5dv3XV3T2XZ4UCXixoK6F6PatLmQGqL/EVEzMy1B2XszSVHf
qhd9IYK9U2/KtNUReQqPrq6u3QrNKnQ1tvjXW2IyjVKebz0zsSfIOaH5q74qhKyn
PkggaSzM5nT6rvP4VazK7XRlOL+flU1sGywF8/AlADHUJiGg1wibRI7eKQZdYB/0
pzDheHZqVw3DoXlsgT35p7QmQG2zzE2potnSkzTC9uGD8zJjpZKwJhtZt792MD97
XMf3SIDSlfz4Jmr2gMtvqRKqMT8uJsJecEmn6UQjzqYciVK3ZY7VKYc2xi8Gybdh
nnnDhoxgWLG0UWCw8EpJRyRK+8CGZOGfmtP1avQ8VVWOpGWc8Mr7pwmhHnD+alw+
+AM2xCjjpfVmO8TIWQHdlUkFXq3l/nti7VNGwF6rv+xyH94zXiMAJonAYBM+WmXs
hfOgkmjanFDjPmlSuhLS6hCi1EhS0BrjXREWo2fWpStw6O865qpYgMhkopDCCsQX
Kd1VjFwJ7kbgS1w4U0rxpaMNK/eLtXOm1366JYNXn6Pa4W+gjzLk+f1R/c24hedK
lnvVCAHk72/pzZ7nRRIX5quUGA0jBHgnj1UlUNrE4dqnEP1jfWJ8gjBII0HI7ywd
uMV5A6FYHovEdEB/wSrkq0Dg4+ptKaw16J2IfU/GAI5G26d1CDVfYITFf4GgWfBv
qfn+Fm7rj8vOmZZtt38RrtHlsCIBRp3iEqJcOr20kaSoZgd4rVS5TfFn78cNRhBZ
1cQhWzOZh89l4SFS5J/cor/rNzv6NIVeD/RzulcNnctWPEuArcNXudWjRL27TkTK
ADMElH5UOBZ+2kzBOoi0vHgRjjwIISBHnz5VKyP2xBEjL5EvwuwtHlmnPZfJ3hAt
3s1jWoVvrMnGq2onWUkWrCM4VEzU6FEyXuTmwurXfiVZWF1BZWyMSyEShtwW1n54
k49MK81vPjJSxAjFDHSttQf6qPDHGGXCE33dMSJ5BIn4akSUPT3RRi5fyEWWiTYU
GBYsf0ThtBwR53z28CEPgyvnnKO2JopLKQ+bVPjhnn0xjTz8Kj+eWxea0p56p7bB
s8dOrFsGe5SGlJZzuiJVu3SI9bsTU2JX6gufkmwtBUxYAMOuzFIqqTEikAr91zfC
hTqOcK2t61J6/4qr1W3mQOIqvqlStG1blEh8Sg1ogVdQCgnO0Y1MnvuAZGwU2lQt
8hCmR8KOOBRcLS02GHv941cl8a0n9QlOWMf30TS3dpw5V29V8jnz/QqrWPZOYvfS
YtvPDT4TzqXiy4NFQVk2QicJlQPdDooFwvMmscWhCWhg1LcpWMwrF74K7e2aIJtS
f6xOdfSaLJeWc7YK8cBSHQFjJodFYyLDj9yxEHdbwo67azDMIZjlabTpSzJfDSnt
9qX68h2AJJS1AUaLDNwdc6pc0vIGXw6DK4ATnkreKfXuYNxc40OsZnHEfxwieX8G
EB5X26O9kcnhD4uR9HBhWijto+KGwL6pNMR3bR1BrjdTRANhfAgUC1EYj7wxboJ4
m6tQ7OxhjTpH/6QKGtCb4Y8cQp+acnM8LlmDB5UqNA40xqxz63qWJWbE10TAcr1g
9h5NNugatfr/jzQtNalHPIzmtgmIrTX6azgOpUKLZh3ZItQcFnXyUaUN+9S+ff9B
qD5sq+LkkOTRKU/l2XdAqTo3RCjmrm74KztWXY2jg+yaXSXsdTVbb93s/6uFkECJ
sNV9F3JIFpL/Zmz9Y1MR9B6KrzoEvVdHVJjHq0Gkiigz+83j9rwWn0+IMFGbBAlh
QxfZ6cp4lEp5W1P/AdjAuwUIrZt8biU5GpWR4xFKQE1dRoU7XdTULV0qalW0f9uR
GgZxinrr5/CCmnhBcJY1p0vnnfk5Pbh152hmLrrbgUp8x4aaDvqzsidipFtFHgZT
XJ+7vKnaUtipBOnGsrFU5gxtgdT3h1NJseGdGBW9/7CJ4SzIZXtz0dCuxDsGF2Tv
8k0lemcOlQrZDdVB9dXDjhEU7lfwc38R3CnQLflHUjACn0YvbXmlLpu4kzlpQWYD
drVqZEo6fH4NBGaGOp8qReess5z3tssDh2A58Uc9I7WWLjS5IUjATPlNxBtATl/i
rgzcqn1vu02nOOxtqfCZJNGTQcpVFNklnKwzhGkJoha8KHyiHBd8xGJWtPiuTsdX
ST3Z/hot+uXVwcNa3MAPlm1msnNcPn56XvRDTQ0SyNJzuV+6lus3X/HGejWaZgIF
RVG7O2drEkkOhfCfIgzxmFXw7/V6eG6IrW2PdOgOdT5+aCeVgSw7/LT1lRXEEKK2
iCwHgwwInODms3Jt3es+nk1C5hwQJwb/dltEwRaLb0UC/AfRy9Uy+OLOm07LvKyE
0CDEW7RvuNxAe3jWqY6IN2Iq7QJS2xx/rn0sszB2VkpNobhD0JOvEIGZjOCnki6P
VP0uw8mNxz44O0FHYQlZKtbuyGR2oTo3LmC0F/sigI8TzWYrivg6iwRHkqI57QvI
/qTnJUP9lJfsyKjx0UIXiWNTB/2JiUw0iAarNRoQelPcMxebAJiYET/HGinZhWZG
54bP60hzAlzoDrb19kXrJzGpU12zalOmU18wXkAfosW7hziSYP+Ws2EUGAOWliZ3
xuOTknvjixM0JnRKgREGkbbIvWMW58LN8aA7aqgibuBw8xbSVE6gFi3qaNBOFaj2
sCZn3j94ejCfacrQXvzvKS2qae9uFJrseYfyTgOddZQMGcKyIHsrV5U5ulckCGJV
Ud/Sl7WSd4SHlXLXRGqhEFF+5DSNLrqBkekLqF2TeoJw3INpV0iDdVXUtA7NYb1W
y2GWTPZpswfvKnQFoOJzCqzhFw4+Ee9chz+J+fomRHKDqLe8MrTNY5t3Tzhm2OCA
1FAt4dPpMlzxIXE/e/KYulBzx4JnVaQbzdYDZa3ond2Tft7EPT2JB9V9WXkPiDTm
D+iIY6LAJlS6jaCvya86engX3j5aCUwJVsatszk8HKx2l0HY1uZP5ezDMMh02NQg
XJJ1XSQOtLgXeT177Y3bBR26YgM2Rr3xCewQADqNVhOJwiZkMvWyWRT7b6gfCM1S
IYYkFHQGVEwfD6M0mWQ2TMKCPnArV27lKk6dxAEFER5qLaU+mSbpcnRqGMjOk7fi
qSGtbbWJggE8tno3VfL+CJz/fu37fkVSXFtomn2+A9yYmnKdrzTxd+UX2F0mgx6n
kFSmgE38mHvr2PXN6uXCI9cW25u/xm0y7Vzj57hoI6NKQcj9YZkPy7t5b7w2sPNO
rQqtEU0W/fb9ryN8ZtPUUcGy9zcHP851+ilo1BxsQ1XPs12GWtc2pLqsNLnlkHMl
vD0onAU4mNuAdZmU9Z7MNNdP5uv00PKPAOerxQ7Lx+wGQDrxu3sSYvvTas2/hu2I
uH+x3pfZCmF9vHdO0aRMiRAZzD55j560DG1HT9YjPsk8cTIiMcnhQSUVBUuTsc5J
ADVWLwIFHJs4BJHyLdhrYm/HCcidOsfsjsDmmuCQA/Jkty1plFiax1tv825RHHMH
vqOb82Jd/hpembO1x4deJUmL+ZGuzMYKH1LBamvfQDHpfxFhIrHKGObwIL4zXiEh
Ppgk6d7Mvp9AttvhdQsxTIwa0j4mi6mFrdXbSTOsQByd9Fv3gAr7E+IcV3bcS43l
whBS9xhN9woRXIE0BuS382uEYQKuDn/zruxQvYlnpWDhmjAU6YqIFr1rlgdq/YuI
3oOpNcMp14fM3XPPSKRekYvp4U6aOccVI1bJt2zkw5nYhXO9ORsY1QTgrGJsQ3E8
lhALeT5W8XSlv5nk1paxHGKGYo5MTsWu0gLfnVrl9TgcX5IwHCRpUxUMSEySglWK
oU6eDDalBCVf4t7HVU7YLUVf5FQp1qWQeTw6ASSWy0H2UsBetGfsJ1O218QYHyG+
vlQwb9KB9tDdkoIWOVauRE0vifb3K9puMlv76XZbKYcVI6iKc3y3IoPWKRQq5HYb
X8mYVn3W9xp7/bpV+TJs9x4FX3Kt/1kRWl0l4VUIrc5B/PdmOocSWNhWcjvlra3C
9oaETJSH4X75RmcjASz+YPYjXUPQ7Mu8LsbtRVskx3wURdSiqvOmClpcHcmy0k1A
cc1oW3E4pxdT4O/5Z4xarkgrrZiBR14DnBg9ARv06Whbc3YDnw3CgXEB47N/9c3+
48vLRYRKsj1fp3hKmWFkSfsGFab258xUzpuS0TbZO4vtppHsbh1So60PZcM00L2u
nWOW2LdiqVx1Cp2c+Mrn88jJZPlxOe/Qfq8kUYVfBS+dEXwYSJgou8wCJ4wv7Thl
BdZcqlch50IqFTHRZ2c9kmvOu7q9Qv+TLVRXuV/Uru5uZ4gofk9JPS6HesIJCaCc
LkLaALFDPKBy1D4st5V671q9N8KgONXAxuasLTfeHLUzIzHg5sawAqTI0d6uGtdJ
DSMAY3Jg48l37yeBdRoULTaTWo3sMiqmwYGXtT5tNOLVuaiEqVrQJ0Rif1Sljqcv
EMNXjHglQtigf8NQ7Gc5QudOpYfSaw57/9+x3v/6Tf9qd3Ov263zvqyOg5sCa0xR
pI0XFsHwvBspxakoirsc0ERp83L6Seoi24t5Zq1zeaVKgh/vRLw+f1UjYcl/8Y69
M8+iDX98/qa9pWUfHo5cjGaQ1puUd6RJPsD26hbVCWqtdhyyBTuRnhsbgIlcouat
paqm/IgXJEGiXPBkDIG57oY26sb34buTGa/nUu6GXnkBbOusu9lHQ+88OPgnjVNz
/JQ1b2FYCyG7CTnRdXlKJ+CA4dN1dlTkDGRNPq5EK/5et+383epCpig2HBDTpA6N
t9YZwnWwm9JHv4u+YLpLT+zjT9M18vstD95zGqRMalA/AHWT+FTT3SzG0Dws9Fg5
Hfk6KRQsuekzHOctPh1SbPBZ3NoIyyN/wCSRaQnD088=
`pragma protect end_protected
