-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ipT/liymTQxd5mQV4GwZIFlbj5QgtrtxlVnkgRsSZ31IpoM+Y4fuqUGOD0w6B7CufmFZvbOCYAOk
UYcxwFuH/9ThxyVWUO3TMIuVyUTmc6NohxBGC8DcdisNZCphBf7maThf8PtD44zU6ZYXZ6xurd/U
eKYudSeTWdqHKkXdR6rPHxfb4tXyt4n2zH2mcrosyn9pMXrCZzaCQoID5TrTzrHbPKhECU6emby6
gucUGAipvcyVyze9moRp8FAEwpNONg2onWTEZ9VCphCXXaE8yw0TaFblAezDRP8AZnnXUg6hDqib
ppmurySpbGOC00BKa0LNjgmTe9BHCBeCxRl1Ow==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8560)
`protect data_block
bLKUR2/oq8Kd7vhCl54tGmvM2GLqE7bfIsp2XfcbS8aY1eji739YIi09BO8UayHOghmNap58CVyu
aGEHnrWANnN1dYV9+50Z1d07lOgCPIBIPN+mHv4uk4H6nvHEVxX3dlT7nm3lZRcCuEkCd1DQbuq0
tsZvr/Ljhbi9/Gf0ofbZA5++Zhb6Aa5g7CpoxoyXE2y3cFOpZEJBYrQG6d04PFGr5zhwei7zpctg
Wy3rQkgwZICRdS3mmXmZHc2l60OPiBUdKxiAbyNEJjEzRo3I2uVT0yGis1c5FxMOJ62usRGf87nI
XPbeYrHcBfUZ6184ds54Teu2q0vckonk1cs3WTKgwlOP6ad5aldV6PppLdNAMGcjbPtIcqO4o8Xw
vhj5+NYZ939BUSzkJGuMysN+2IN3d6QQSDQ6nSPhaOpPFGxPlVYO8REHoblyV13kcE/OxzYUXvnr
G55nrkNTm1oP4At9YewP+QYSdB6CnQXG+BxFDblh4SwVsqZmse0fL7nFsqGNvAiSbWGqRwJnT4HE
GQ4byVHD7nP0fhbJgoGWzpEw+OoFaERkaThVUVv+IJc9HbuWaeFKKjrpaELoL8o1OaIEKGwC8hHQ
UajZTuMdH8RNxg2a0WwTZYw4ZjBoCQLutbLdfRsj5RP3/CdAUnMorQ6K35whOtUSltL64RtJpsfD
3cNPROveTtiF6NeWnBW2oGIVVnNEKPS13x3EyeBzPNhUI6msWAqKvgIMiLr0UokQ4XV6qAh//y5h
90vE07wfsN3zQE2LbGQUebj7MBeVKaSUxcaQM5ieoATInhIAb+OcEFMvCUl3GMPdnaoyfZG4kFxk
JZpxGox4g8FhWzKPytucZb0k3eDc+vJ1kpaCT1NqyibWFR9fzPDsyZ5hTV5xQDAlM0F36sTzSpFb
cxrcMvoY0IlKeFGkhztsjv9DFn8iHcogkn0ulY77SezACqmCGY2mOpXeCSN89etYbydThPIm0DoY
aH7q66WjfIWCxpdrbJrEwcoAnjyr/hns3YhXo86mLmXpEfxHP+kuWyUKUJU51VRBx9xZHgx72758
JNTGpJRCup28x7O45w30NI7mQ2koVOWgJUOJD4DXttfNOzRndFeH1uAC6FEY6WCefqqmjBRBkAHS
yrzWrAlFXoMrVomIffpRjY4WC1PysnwB4OUz2/F7aYULOA0HTQzk4H8ImrToBfl9G3sdXBmWRq6o
LYO6/MjDLOPxB2IqW8tCaLw7eWJHp7ruSuyvbUTA+lVmyIsBIOuAHiSh628YyUgMmOW2yhUTh1DQ
V/EXcRWuphq3szqM8meQuppdUqGC6jGU9KSFMWcmF9vi+iy1/JfwehVLk7Wng8umQD8EKwS654HO
s+Gya45UdCURyjAEeuKkn6jCXy//+2Wi7U2Hy8xTfd6YseigHCBfrf9QvbstFVrNcUp0EVPAunl3
ZHwhIn1MJ7kKQLGSL0v96OBcOZxSjjKGCvbT0JhaShLcSagjgFvYxm+TLmyIUp7YpKteMoSBHJv4
DW6nvOyvvoDwS1yLcWP+Agj7UAf+GnGpi29iwA1OjnROsy05dCwHh1mww06LCifRcSneHcl3yfSG
aJqpd0h3GqoNy6Se5gPGeMYs+pCERhuMSVg25a4jePR+QSvOZluNvS0coviCiPvi+3davBgjagkY
2y51f1YbIL8VEL2s9cR6zIZ+yikOmArqB9LlNhREH7rwqlwp8QtYgrnfQFwuCWVt517kzPdTPHml
MTmcr5KSiGoNaiwVgpFJG34EylyaYRFjPHH1RK9Wa3L1S8/lZ2RXe/TAA1vxMpKr3G2PJC7zUzsL
984i0ftphYupmEGLEjhcnmYg+IvmxqV+xTwcmD9fs3YyCZx2c+NEOk090WcfiCl1rlSOXxO4WSbh
J44j7sL4uAx1BHtfoSQE7woCxfkOUAVPSVjK8x8dDOMy7A3JBbe+6at3q56zzVpfQ8ggEXu7XfFO
J2kI3L13CcHB3K12dharzqF/DPgEUWCJOA5dPOqQtkvrt1ucICCFHDBaQEBA8CXxpBxky76Ig/Wk
MutpCCPQlKMnzMyrf0EqzeemsGUT2hCblVs1D07T8jpM+0e7rS/HWiTzznkvEoSvNlATCUG3nJVj
efFe5QiA1yb41faGCQayLVdl63A6yhba3r0TRXsKBzxvhqYSMtLkThCflnf3rLe6Gi7qFcsTBMLd
11eVx6qz8rcJbG0uy75ll1FLirNgkLFHXE1tuiTahpuvm6LzPnEFhyCyI/G/LkTfHIyXLk84uWwP
q3YYqWedsz8oAtgYhKNhYHqKiLjgsy4v9dE/WNVsGGJMRjS2zX5f2WbKcp9y4l9Cj5reQwi4s7Mj
TT+Ql6QskZhTQhzqYe5XslrsMBK+aTNVcupzQQiVsDa2DwITHY+S45RKbrG6XinT8RYVSHIRZBWZ
+MpfAWkJZtN5BdfhExPQNdZ8BMFO5eCqiyS64l2t19i5c1EBgqpRU8kuttFWJnbfWpJZfrPu/RPS
MoNQ/FxkOlda5Dyj/juW8mdEo3nk5jJ3IrqLmnW6pkw92yi4rZ5qRd3tvyT4YsCMZ2vXOUSssGU7
IdImyE+5icoyGnLyglQeNZlFjqUkiLGkz9RBJoIOGYLIcpTqUEyGUTHW28+zxzKuUje6T4IGWQcS
4mU0I/z+wgFa+0RtYBQjCvivGZoXCNrUgq4bNUKn7C74BI72Wx+zPZtY/fRteqCVDicqQGXgBFJ9
G0QRYE+IyEKDMbGoqO29Js4t33yjHAPdkxNJLoEKOZATmLnuk0aIopepF3U9AcJLIc8awO47gv7W
77updeBMg39VaXmN5JClWBj59hIZkQV52O21VBFOz6E1LWwgy5+PGM+nnCd5OMKsWY0WUnJgkEgR
6Xsium8pE7KyDvwJOo7e6NrRN/4zMlRaUD8HL51zMVj0CIap3XEGZwJwP9Bqr7x1E6aiEM7Fc5ge
n4mu0OI1PwXN0gZRcghyYhm3vaGDvtAI+LQ3kcosoMM+zwkB3oZ92BblkK/ZRa2rEJfck7wx+llX
HvsR6m+mM1hbiaEfnY9I9k86qzIT7OqKPRbo4jiMw6/Q1+nyNt4upUek5oUonvJfBr3QgZ2aIM/n
lfQvhPURuGDVBd7atFiRBJB/PpZElwgk+071ptOJpRdrUxoAyOji+OQEoRCkZh6ARq9spg+axhhq
QR6Dib/xKrgQtKJb2p0r4uuarm5zQ2Q7qvA7KdT/0kL+bZH0nFmjB8WFNk3MqpSAdHdH+CYSbQU2
MFnnW+WMMSW2jU+7RPZW2bqKfaM6Kx+AYE+RvsAImP2n+0UYGracFvmZ0H1RerkI1/leYRPgW3c5
vrc7zbjLm23CJhCUbZKx+0DEHbEbSLXiWzF+D29wlND+6BKqmndDWA8hhMAiiwuFJkRYD63m3Fc5
GFW+Ldy3tSU5GAx7Ll/b9TpTj4ebn5I7tVFsLR/RQymfex1Rwq4/bu+5Qyw8asARbJAAuXZnhdqn
lLONFmZ3wxdthm1GLrIShikWli2zm+g4GBCZeW9yfuRDYEw6QfmKcXz/mU+y0VARvYoBkulTgnXR
L8uFUqQ6U8bhB2288A88d3fMs/1/fCFIIPI8Hij95DYMJJMrCmbuVsnnP2g2AnqMr78Ib1qkTxjr
f/0oMZrasrCJE3KNrXd9iBLRlHboofwEyVo6lXuH3SSyXeJQvq+PYZPJtM6ztfU3+BkkodsKDgoy
UL7aESqNQI3HTcK5oC/cVOVAni401r4KW2gVq1xBeWwuI4WKKvwEWBvEGxTszDlthCLCtfLG6yU5
/2j/Eb2gD/STKmBRc4fWshM3lZmJmumNh30xF3uMhd7BNBjdpY3bQHnuWQ8r5zlnzwwIeYYrZlOc
huOdz4C1/SCkwhBeW/7fdgU+z74Dt58EScbOiHcC9tqVtZEMku77avr3NFNeaxwhAU1BfS0/u1fu
fkwnWhDhDPiIWMDQ21rvTjKOLBX3aQOlHlJqrrn7gNhG0r1YPFgU7mp0qTotHS/OuMvhglhM/b+M
NkPTLHCHMMMZvDYt02/tgGvOuMZjOuxRsfNjzptt/i7iOOncSqJizEXfewxXsjmn3D+leVbeY8nu
O4QP4KXlPiUO8XLRAyS3D/HL2Gydvjx6DXVw029VojVTkCT7nL/VpwbdYgkG6C9s1Qjy47r1VOhr
8j/2Mi4DF6AML6lo6Gt3S6cjEa3ie3OoG6eOego92GciH6V8ZuJE1x0MERqiQdgU8Ny3X3Yh82Sk
Ly96NUoRRigxyiitRlUR56dL1JGom8QIBmqviq5O5ijNsMwYrUd/tmLNDynyRSiwm3syG6gS7WLF
DmHSzf6LV78a2eh+zHLEjJwGePQgIZBR+IArGzC3QATCuUl9CTp1QgdvlpB5ihAJtSV6ECz8PCLH
CLItJuqlnJAnhCvDhWe3bczpDRyYtQ3o2kLwDKIS1AzGj6HKMywujEeGgqNQZSoIVVHR2GEkJz58
Rnvy+EnkKydePMbiboIBKNPyLMggijzXYp4Y89wnA6N0WSOXZjwtymAeqGBEOSQQplux8LwOzk9y
Qdyl9Rjkwsz6O7SxZb6HoN43dQgmqo0VTMI8OHcaxC9G90fArfbIQObti3Lx38mFiZcvZFC2yZm0
cD0DaunnfOG9fX+XKhpvSotrFV81vLxVoGdVyHqhE3+mDtDtv4lZUmuYhDR3/LUduHt9UDHGoRi9
t5wB7VZHiHJZ7VdGIWgrLWjxT0EHXTz/ZQ6zLY3iUl6xz3lrObSugjRg1R+YmbbB4QzYPIFsphmX
GKjrdVS0jXFZVXN7TvohjumlhKuV5TUkeJdoO9gDr9QTbr8qjH1hIlzrCUDQqaccxjrY/NBOMwNR
Mkm6DfxtUYvjyc5w4MuS+eQaEq0syY3Bdl92F+DABwIfowWE7/mMVb+cUTzaY7kDGDvSPT6FkN0/
jpN7GfK6xQqW2d2w0NOQGDlfq5YD2JfL/XdSOBVpIc2pfIVcNOPjDOLk2GO26Z8xOsyflriel6d0
jvjp5lIrNvXtQ7HIVOeN09xtCPPKryrPPXsT2b1VV8cymepjVBViHsyIY8H2Vdz6fAJ/JDgbedkM
VyqPd/BJmqsA6EZlTVaXVUinEGvQZTc2xnwVBq6uAiaykleR9dXQfTgG1eE3KfA4FuQIvcdIlc+q
uOkDDOWInUuE1zaYb1mjsCVDzevlimsNV1Wl9+OQF08FUxhp1gHuj8LtoK9an/JhzCgrhocZ6gvt
U4aur0W4cWIO9lafREIy8EdTF8FjyjvUy8kJlKo49Z4JT5uBeNPu8RSr4zSlQLKPBvtxORm+ngS4
Zl6LnLd9cym3aULuDwWmsGIZULVSEYe9K945IV08KXa1ASdyxa+Xi3JCXQFZJqpjFN1j26PeyjgH
w21V6hlTqe1DSNjYCA2A+Vyjw8onYTFX9niLaYFkNnElu8+SrSUKlhhw9WNf0CENDdvF2BOMyY/R
xMWfjpvdJnEmL9V5cLXJXNhSpfk1SnNdu40U2SN7/nKhgzVJrr5+HcE8DpCPdwD5iSdtIrvvmJdm
VTK+fZoNUIDpmQ3wEwbSHblRfSbFn6JVb0n2OJPPbBNCgh09D43udELetDubPpAq88RIjxEzbZbg
aYa5hPk8tx4d1q2O8EFBz5DDgqjwxX89e+fh3w9/JO13UuI6GrnWM7j5bO0B11gVqYeqOVHw6k8b
16r1SYDx3647MhT7ZY4Xk1+4m1gBg9BAfGzKggB7sg9urBruoN0RVAg0Zx0KSATkU/3/IpzxaH6Q
wzrYXF5N876bhASvvr0/+V0/MuHE18lCUedhQOOBSp/wf3jtPY+MI0A58gAwiSDIpASp7j6lh0fe
VIH+Iiur3v6y5vs05nYDA/ux+ytysNWxwVlGO/tfN7qjFJskLQtb5bQK2my6soKwbuhNlmmTg+FI
28EEGLcHiqaAADsdKlXnaFBN58McZG5Mv65eBhhvkS0xgB3verES1f/r9hgcdJWDOxA3rbmCLveN
WgjpcPFsGYNsu9mihDuhYV9xtoxLoH8Qwty11ZS8Xw7APDrHlwtJwhCdeLkL8G4654/h7iHKYmT1
HVCsZiNy0Z2o20sEpZ5C6YG5KVDRJliu0+cmlO5S6epG400ZcAUxoVHZY8xDpYfcmqjVXXmD0ky/
rdDf93A/vVHO477ktN4WKtsX0fHPpkcmuxWGf/F1pIMRoItmGOcKeSoo617DVIsiMcwVEGb0xIb9
j336Ur3j6re8SQ44purSiANPC1V9dhRwTwL01rsy6Uxr+D2hv0JgVgZnH5rr4Yk/m5+VVVTOAL6b
Umpba8iLbl9HCo5ihIBS9fDq6887AN4ObgNekTYUXA8yJS5+6wyHzenhATEUJn/Dm7hGquRsgvWX
KS4ErUISo/MVgEd3L8vL2yx2Xw9eQCc3taTdqaQUsa4J38btk7MM3xQZ4KMc0rY26JyqKMZAdVNW
QALwZoFhrExuprfYiVgcvu3dRkiG5isMr/DjcdsogXqPdsrSGtIVaOOepTDY3KxrZaNiW58ArpEY
9DcInpEmAO86PvJAQ5wGt1deL5MvL5o+4jIHKdK3E7CaMy+xqxNq1b4HMk1FmsXJ3/URiCfjqloL
GvmIpaZK3rHhPvifXcxcloZxuexcU1snvYZcDnNyXwQqMK7fj5JH58QxtkJh8n+yx5QUs69xPE0W
/bYZ+OxsUZkL+TLJdbtxB7d5D7mhV9GdB0yyTJ0CWoPisvJTIkLsqR0i/ooy9M6b35f2sdURwuk9
9Pg2/3suRBps1urJixqaLlxOFVdPt2srAIX5WZ5fm2HV/9yW3jjhhOiVDld5A98ezoB+qsMUv+6X
wBX99jm+Gz0pvhMtm1aTSl/z6uEjz73y/WiixUvDQjA2W4l/1KIW0dqXSJVLzGyfz8tPUNZmcIni
OB0Nb/FhVZ714HK6aZBcDuw/1tT5jw2KAuBNV3F0raN+boEk2AJmNnxnTH71g0YKd+O5Cw3idH1U
cWSlsYtJ4x8h0TLESGWabCn3llq91zwvbqklG12QAs/OI0/gS1KlsWIjvE+OfO564uDFsezfE5+Z
y6qZsALkqMtwCmm0+d8vdSuT8hBffXSrhbiA65lvDpSvBdmiZ/yJbGM36dGS5RO5qRpCHjQBK8g8
hx7pjuFibQ7lycv2k83azCHHJO5gfW8yPrq+yBAqGfy4TsJdpIvha4HCFkVRm+eV37zXoJgwQQIg
TO2R2+FPcQoa3wjq+TKk3wUuI/o169p1juUSKloD+3nxOoPybTn2+3K8Xylah5wgsarIwzhI+GpX
sk+crnfLqk32shBpg5kT2TsdGZKA6fS9jCn6NzKBQ3qUBt5b9Y8kWqAEZ1sRZgHZ5PzLveM7p/Qa
YHNni+QcZXiZHaR29ruMj8BCyqGn98kuXaq7OTewulfJ4Hp2c+jnbMwWFWY4dHUXslIY6rzELytD
8zG3/m/f2aojm6y5xISGbZijZcPTuX0jYz/6IQymIAdUrk3zatpZVqlpgabLWw5le+Ydy27kNGgK
TsAcM4G4daevueXSPp8rQz6Lw66UR1DJ79Jf9HopVRdtPFRD/hYfKrRZhDH3D0hrUky8HegTkz6u
9ohLQh6TyIA9xId3zeyCTXz6gnh2lai712LZoMVLOK6I09bbBwJltqcB/UJjr1NVctxYPj51FREa
yvi5tpYVKB9snfz+UuB5050m3MJNWTGeviahbFK7dO0c4KNCY6KKmZYgPLrWQH1V+3Jbut0LKhlI
cYHXjjYKoW/Q1G0or0oGOckz+2CqlKds3+pQazFQmrDqtcHa6A+6NZV7VWMkoES0zOUG+/WK+1Hb
dH2gkl9hYlPP1nXtDuf2Z4wMXjptJ1r1fxng3DYBWW7tpZXu6orpf/I/2JxiEYgIahuNWPw0mNj5
lvXPI1XMy1Eik93T7AVqIO+2mf5OT+TRmeCGYUFiXoVeLrquI+4T4+HbsTF/oNSMeJwQVF1GgOuL
b8rLyztOQbnYMrid0f08kiz20Voj+7fwm6jreyWg7TOvnxujwpQm1JWjd1M2KhSHc5uQT086G8Zc
5oxYRAWJpkDdMj9ggzldCi6DN6AiiQf0CDCfzXieDR7jjtBNg18hMjdQkSgCbvKNL3EipsAzlfFm
LR5rU15NBySOxg8e8KUh2KMiO2KE5+E0KYTTGUyVyg0VlT62M9XxahRIOih8s5To5n9TmwQA+HMA
hUR97xC4TlUs03aJasaUJvEdMy7lWL+CSO5q/60bJS54L79xPZsQI2qD72mawVz64MwvMmvX/VzX
1TeaFkzeroJmFeGKpJn28ZyD05llfg3v3etCETdzQjPe2pKt+bejW3XPVeEZKrMef93QcSEFDVNL
eqVzbypyAUsVKBk+P6vyY6m9vIJHs4C3Ap+vTLi72+k1g/l7HmX/LHLd9Gh0nZIx51NPLqgZbHDE
79VoyqO6Ls7bw8lronwZLY7669sN4rMsWR3UQpyZKImtDxzxG/o6zwgUwsV8Qqvo3nubdXW49lJB
3b1gVJ95CLvrVvWUs2t5ty6qoJzysIajyvh2Ah4aWXfpc58N+9rc2ok5JR6sADzdkwTcru1oJ7GT
x1xsN4HWL5jWx4zmfPoENhYt5tj6eFVBHEcrK2qp7jRsFuTFbLa1aLJJUAyMsP1ztcjY7nAuj6Ge
l6uXagjCTLx3ownZQBgiwMJ5LgNDlvxCcjSUWwDgwHWNm4G/8HrBDohKK/OFYvOvdwBaQ9VPEyGq
E1zbdv40i3eiHthx3dNeKLHoYw/mtJ8ROgKgzAyApvrdSaXbx10MRPhkWuuVbZcaNHRy2anHD+tm
fN90mHKL1BfmYAZMIXeLIJZn16g2EYUaEWwUMuxd1qefarXF7V/hH4/koMEnVoz+J+v3TcPW6JEm
Axp41XPHA4b2rii+uxrMx74VtFj97WqMEq5Rn1Fi0DMgqDMhjyzxK1/xUCkdKlWjXn0Joc1vtRfe
k7/6Oju6YCjFrMQ+rscpC+LO+vgrUR/FGWfcpcwgivYlCGd1p6chPsPOhoVRpXNp14teTa7130v+
b8J5seReuIatSLitGO7kFZBoOe3dJXZdDQlacEJdrtu4KtJikPwoJYieWHt4watQl2hemWULErtr
JjoXDAMxo4ay5a3XKaq8HqCVCUoBZJd3WUQtyqY8BkOr/6bPNAwI/W9ei2XN5gWfurr4oNf1TrUk
VmxD7Y9W2+LR1l/IB6ditJi0FFNaxvnUQiaVsZNtrFDH8YtI0R03oP8qBZIoq++I5LQrlPp+buZh
6He9RY+QS4krAKXNCodt6DxmRLCuu1WhWvgFgvyHbqFqist/DiG2r8idC/MJhmmyS/DSinzTUcyw
OPi/cP4USoODvOdHHW+QC64kMZzCbbMmJ7/QyoaQfC8JvpVQF4g5pBs5dPjhG2dYuwod9Acb+Di4
Vtum1eYDH60kb0okh12dNZtlt8EO23e6X1t5vHd8iV83P1UpJ+rYCqoIQKnyGotSDLP8zBdpnceh
YRK/I31/wS2jUSHdVCNRDBkIgHELu+ZBu7+7qrtDb85oh8bC0tJMPfAdNQK0Ozc/boM4Q+PKoVKl
mJZdhVs9R+U6wT+YzBwvz6FJOWsADj+W73poXPlltc7fhl7jGnttEkRRA3H6Ihij5g0PO//xhFJb
6GmoGz04SaQoRiarmdNWW9lEHPueZTu2V6C5c9hl6P/xrJl6p/87WxPiHeKeTb+8V2WNI2XrQZuy
wxPwwPHLqpqEDYCHGAd/Z6KOb3176utFRrLXmwSve//Wl16EpTPXFU5zCPYIIVjlta8zpFLqyIa9
LkKtt6BMHrtRvq1R6eVAqMWTIqB7PDDlFNH9JCInEzwF72IdF1N02+oVLEbIQe7QyowDdtSINc38
NdKpy+92SAmKjdT/0tL6NCpxjMsw8Jigj5zFx4jY8UeR9Zds+kGA+jmZswgCC3t9JovXvRceq2Dc
hhWaNn4mZO1Br76+bVivAuzWb8CvpDst1fWSb85NGo1ScCD+Hk25wOQj5zrQ7ncca5MdlC9EbTQn
JOq39W6l0qAoovEBEQT2R1WWjFN2/g48orvKpASuWfqYnm/hCULbOPPhJJJJQFbXFDOXgqxMg77c
Cz+gZan5J/Z2KD//vFu63Vkm06jTtf/bMWbkQqK6XEUuQwH15aK/Uw00tj7F7Urbyy+6WvwyV3iV
xQAavAtlAvKDDD/N1cD6ySFiTCjOaoLkKxihXPorf6NttFhIZ3xk+GV/HAWL/7WZU53Elt8u4MXd
9zlQhmDw6Sxii5vxWePneIA04BQjZEYjNfTQ1PrGrSkH56jZYHe+ckP5XCNMR4ISbFRT0YEGLk92
jv56CilMyTWy/WI/QZI6+MJ/7vviR7jNvI6YWioYXtjaMXMwvDPPDYcyRzbEYU5VP6G9q52sCqss
atQkqdtyCb/7BjrYtJa2+x5XXXDANvJ2SGGhNwabmSLuwXJ1iWEKfVvdue2r2Tk+i6Yc8MItBm/R
97CxUHoIbisTiDmA03l3n15/egb0FZsESSskSYG+O/yi3+Ra9NmxFLOrqPc/ossNzMOxLblcYoE+
MPNze1OFRThjCIEgQw0vUtTBEDFht9kn35I7WrBe+oOAIqWs9yyDoVFgYpr/Qb8SsXPIG5WjUyXZ
ZijbxNthOJYD7czcxPi4v+ZpYqApq7uNZJBNZLBtxvt5kOvUQ35EBl77bYMbuYHgE5KJVe+VOshi
TpSmrSVk1lmU2eq+TvwY+5jkywja2wc2w6HwyIG4jBfE0XM9ASmYwQfG6m7iATrHY1Q2vGgLBK99
kXaRlV3B14VxY6We/XNYnDwF/FeSw5qMxI4wzqp2p6LKGLT5V9YApTOVAdscw5lqaSqjiTwKQuhz
zxcibZi3uxaRnB09m8OBAamXdJLUwThml0l9dptsVHFb8yEJK+Nz61weSYLRnh7xjwK/OLX4CpsP
2R39C0MyvwADAplRt2dqrPtJE9b7b5QBxo9f5FlwvR+yHz92IleLden6tMjjADTjKW2Va+RIeVY3
mHK8sqQJPpe5kUgKLOyU1eG5wcFMW5zY6EYUJMR91QLg8WLVlDB47ImyoCVt9G+OciDmLyKAcX8T
VrUIUx1MTuWfqxDA/yDeUIH6lG+O0XBpM+P8wsdLtjnxtH5GmLhJUANMsFDlpWvioftuIqa/OP3K
CUMOgms+skG+o8WXRgBBRoBJtzp7rHIr2tI7Kd4faKwKqr3+5zLniIRMgmbf+Njd6iVjMJlcWv+H
mH8jvJXexcFUnJ86sLqQg1kfd8btGexwOyXk2XibgMoxTDFoWOupKNU/9wiz7YML3m/vH4Q3d1NI
HKRptRIguuG77zTTxnFZi/USBgKrGjnb619Q6FOgCSxp298Vc5jKlQl0PMeoeqQAF6RpsYJCSvn+
YH9iBRFtJ2Q+xg==
`protect end_protected
