-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QnKFjlogwKQYXbQCPoW4VrpOfpWGB6Bhs7PQbFsUGBTMAgjY6Ao/2JbCk7HyZ+0az2fpYmRVszJw
D9tzEmeVgc4fgj88PrpID6uY4+7AVLVA5ZXQinI6bn/pB1AgKSi6SOe2tDbWKBScaiCiXjGAdycx
Wy8RpzeVUDyNFWYzRU4MRN1wVq24JP/ien98Z9tlXghKtSfK2cXsl1GoJUwSUviBNZPYzDVZwr6p
az0ciG2biMVmqgoyfZRTSwga8XmRVpVq+cwvjZr7PQSO8/PItLWZGVB4KBs6qnSIpWq3ekfSCZSn
oPbXtsKc+0g3r/byCVSghXexUbpjkmJykcuSHg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2640)
`protect data_block
3YDbK3WnXQX3ez60Ui5djDGgdp5KOPjssiXRCzAhqPP0+vTLbVPZd0NZwnxSoWvKqlciRgIrb47C
IkvpkwCnjJnCjp4v9VvSoIt65XI64jcXWrZ2CetiLfZiCUvkQyJ01B0BrYe68gxYXotFFtyWB2fh
t+6zu3PELnGA/pUVe2ssy0aX9p6fGunTquMVe0NKj56l0WbwPGCz9/8sIGGDFZjsj32YQa3J5BaV
VgYZbjMM5C7LpJAZ71zkTB9ZKqknD+D+e4W9nngn5UwnhA+g85dyEmEQvJ5H38k9Dr3i8uk711rn
IgTyqV1SjNDbqm/dhJHxlky4Vu/uGZeKMkf+QBYCtn74CkaeXr7tRvK82zq6u+A6lWeKk+15+X9Z
KMNJ1J7aqHDQb7558xq/99mB03J0vbNhR137qIE5fgKzg2t1BgK4tbvgfv6BMLVFZtIakyFsSPea
liDKQTaXwQXKDoHd1RuaYLEC7L4bQ1zmvTI1jCzCGnfrqhYRWYFzF6f7Fpq6gcQbT982TAnrYQif
Pl1yHaReH5JXjIA2iLd6UlteULEoMd+RTwu7DfXvgi4WZjCt39m82xwTpZmcar9aLFUX3Gvx+7ia
FlJNkBy9EDhXFo7PiryAppvdK2mlOCW+ZAHPl/FAXLq4ajvQRA2jSVdwIJ78LVDNmzNqaSY782TR
NhRwYStk/SVdyeUgFu3K4KQEts5vDY8+Jy5zfgzXI54hYymrRQlblmfrQ7XbnBGnWxDJC286WLEE
vGSKkkTU7OzzGUL/ML+M2t0V1eAv3lHiNQFAve+Ip0rwu9Ci5prHRqs2XsAb9tU9gpz4ER2JVDOK
YyJSQHyLyBfb3sBYK+n/YZN2g5WsgFxU0WNHIHHPCVhFeMfuU0Or/x0ub8CKbFdxj0qhjC62/fi7
2zrZYhlp6jaFR+lN3wwnv3yGl2Nx4C9gEIfHz1fhWX1Hj3fjp5li8biQC9qgxrBHogwQsdoDR6NB
SoK2sEg2a81ETttggUTKc9ChVo2GJD7bNsc3PrhOpcxqkicBOlIRp04Erx+jc/O2DZ/vpV3nzmNc
oaGcfSK1ITOyX96p/v2WysQapmoK5aFRIr38EaUOokv9PlVpjBwWmU6QNkU/5cDNkcr1D9e19+Yv
QMKKSSJWAOO0OB2RBvq2Zu6+epFaREyUOE8PDVBo9Xd0PS58cKaItMMGyQp7P2dhrV5IDmCXVVjV
QdHBMGG4l8qqiFBis7Ihbi9lSDkH0CJE1mlb0W0T5WNcJO2cK35wvUzSG0k7Q5uxbzO8sp8aTJdl
TVVUnFn64CSRkgq/LQyaQrZF5FKyxIxP8HGrg98BDwsMZ8tfmG4W6I6QWAo2SiFheaIcLBNiyyUi
KbC23+13ixKKC5EG4ocL2uWRfY+gm38VkSgJKQ/XsoYzTQEWTXdxfVXFdasIYyZDoLmquvWO0OjE
HhLZk4x9v91h1wBAH4BNxJGftzVpYiOxrG+2tzsSfny4W+Wmf6Eg5WES8PiKS9mPwnkmTuMhwV38
P0Hh66FAtZRCp8dX57VAxzkkCbi1bzkUacgOGgYZOE1q3CuA3Mbg980tUvrNvanG9dJHU6mYilNj
+p2FuC6JE4lAOMNeQdVz5zlNxC7NVJZDsJnDpUj0rTeGoVwYCfMlMn2Go/tljPMNRnU9FYJgsjno
3mnoV5OUi9g/sNEooxQ74Z4iSS5/zLpI2pac3BTjWyzPE4XKUH/9nUlRYxm3p4VgGbwcYCjT9nOT
9h2Wx3Bzg4+IGZMr7HkEO2NwFX0eoDaHZTSLgpFGPoi6uvAWCc3QTTf4ZuGcNhzoxonpl4o33dba
pjum9+lEau+mYglyB9LWlHTXv6UTjeu4K8NrzwPh5RwxwNWfJ53q+pjSkwtrYIovP+0FRrZmOH7r
/iLI2r5Z2oLMmXWn/fF9M5kE0LB3JdgNtOQ+126cMKDroWlZ16yCbY7VSGwnqWI1FZaDIUUGWcrd
im+rKD9Q1lFUpqBY4RvXsTZY6zQLXGQlPRDTI1vXW096NBJF1vJ1uGRqf2vYqR3LmFYszzR6uUm7
pvPdkltIswEy/ZZNFspKADoLAL19GylirEi96Zfp2Y0nYrhNnuVJ80dMAtoD26cRH1yTPSeWijnD
s93cd+lLl/qni16ZJxN+9cFGA2M/Bsym6OxEjkQNKivFJG0p36byJk3PKOvNPMxQB3eg0dCvZ7gm
6bAsNkyYivRCx+lU7Yi4YWRqNrBs4x6wAQt3n9eM7i0pXA6CZCgfQdEhkZpF7QdCwKb8YRh8d5Bu
VjZQa4QNEMbm7odkWoOHNpYGG8FG+g0gi3NgjPsN3XupY/mC5Bk8mFU4+kcXCUKxgx3V7cYxiSs5
GvgOw/VjeUFwbwvx3mTLV+EHyYFpg3g4nOU6g+u5g4BFeTI3wMHZNOiz9lVgN15EPt0OS+s3Az6y
aD2a+HJOE178JKZrH8s1jcUcX21cnJcKOZqrmCcC6os3UmZtC0Th/6xu568Uz20furN/Ngx7mrf8
JqYpCfNbTQiqi0nV7/AZo+WRPmc4CqpsHbPJa5lhVEIzdBeSafXp5+SREdorTw0ckAiVbTBJA4mI
4csLn1xsafqnUbtxE8+L+eiy5sFUrgz7QbbfwXW034AwKddnuUC2Pf5/hR1b0z0XURzJU2qoYOsT
p2ZQlzC7TV/St856MrEbzl401//1i78PqStRjLgyWn3A4WKF5WFTd+UTllnSoUnFa1fWzVaxasro
pAiNyvfIaTyikiF7S/3nZCuU7B4NrdktknQEOtKSay2Qo4a5MF7Xsi5TfQJV1Ul4dynqUmtIO38Q
UNyYuY6/pf+HME9GBk3t3UUArIiMfUJyY1TqKT/vjCscaIlTVWAMJ4lC9MvvQSCVdf8j9cebFiPP
70S5T0/R+1MnknBf7T/dfzdwfMb+6r6YXII3s4uiThF8Q4Zgsx4GvwCWL90u1ayG4l2X2i0Armsw
Zq5W3hrpYlWyHfgCDDefI0MMK+bDVZkzPo2yWHcCfqf60R82M3PsR8C+MljgSXK7CYmvChgxNNtJ
wWkS1SwhyYHAPzmcluyDQCSntjUPahMa+dWtlmoFXD0DkrkcUyZXGB163sxGIeq3KvzrdCXO7skD
3QfrNgyj58d7OqQ39AgfZ9SN3d8IZ/eDnoKDnSx2V8qpZzn4FGX5s8fi5VOoHHi/JYjaIDnq6ko0
IX81M7H1UtFXGuGSpPn/q0kqtNQPsHEYi6KsNGlSrttnd0Dg2tHDhHHZTJX/wFEKlrYSvcizLGVz
4XqL9EzPMXD/ACZFjSWSh5yBfncqc0lRN9eUQbAt2Chd2zrLHCy2GNiM/PmhWqlIGN5exLZd67h1
JZXVOiEu6ul0Ca8n/fL2Hbqe8Fn5KHO4L96CcUmRaebBvyJQM3d1HOjxpdFRl39+4WKVLe6xdksH
VMJrdli71W69O4L4b8s8/w1XmfX1sMeSzeeojwCBRMoyPWs8Eg9lkingCuWJa55LAeUuVE5L+J00
BIMiWjNm9X1RZ+xB+gRLbN1B
`protect end_protected
