// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
AXlsmGLqvvKYHmaeQ3OARfcbWDEon5de3K0YNyxNqFwG6vo6XHhHagJC32VFpbzppsObTBHXvFpd
WzxXGThoITDE/x5aFUezDwJNwqoaXXMp386QohY7dY9enBakFpZC1xucuL/h6Ide9kV1MT5FxR1v
uhCKGwGDaGo1uIWGBnVwEB40kTBrtq+T/CxmP1Ozu6vsVKAp2rtxsQy9MaLI211YnChSB/q4KkWG
DJXKYAFdYxTIH+lPu5EExO+v9mmbJfUI9DCR/Wb2+K+wHpLkEF3CITiMu0beio5oUaENAVQWir3m
Tnuv/ymMG08FKUCX/rcmSE8DNR1BKk3qIPQlFA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 1984)
jx02E+vL/1DuM43ZwMJJzxtcyjMBXFO6rHeIX2sCcs0ydIPT2h5e+iDoK79XJf/ZH5N4x1QRwvFD
YAIH+Rm5XJrjrxztCrOWDMeS5mjo4eWE7V6JPpzzZdWFlbTOYhQnXnTV2WYSQYH1+fI9aBypvfC4
1WwjpHzUQ1F+OgVstC0ut1vDfdBEjlNmAATvLbu9m1/112nmuhtomrC24pYoA0Io1W5WobYdjmbh
B6qlrS/bMjSmNuIZ+HaIqjSBgKzkMS2I4yYHGHsfVg0V4VWdKUyL05x1diGiuYjMUhZU8n7KiGQs
cvF8c8WrhpPDZ5pYd3vVg/vPuJI8NLtffcxJO8eyGh0/pUEmQtujaGxuL4+8O0xn4MHl3I3mmkqr
nB/TvKmFu3bO4+oKYi1Bjg4hPBzhBCvO5bqX7TbXrmNj80ADg/SgJEPUteqSxDZfsNQH4bKh+dfU
LNiqL1FfbN64D3Ji4uNES4+E32XpY8jhYEpOUKm+aKKD4SwBzK9epuwMm6LXbXIi9UaCCA60un/Y
fSPLWmxg/SJZlFIXHpQceR4YQEvXvtnk+zhDdyzSQtjBOw4gUBE2+qxGmjSIj4oZnmPTJnJsEkGQ
r27ob/9QcFviWs/MJo8UxCafoIM+3/ItwFMM2EyvrAc0fNq66nyzFGThGtBirhhOQRzr1h+IknQe
bQsAXuQiVNXlOtSKEN8Pc92xYsx+idoMOKrQK6Iy6ON4RkezydzPCSt03z3jJyP9V2Ljset/a8J9
nyzFEyF54skymBLSvcTXrIF88D7dJa05u2EhvpfzkJ3e3Jnt2huoCXXgZIauCsXPZyXVt0J0J6z6
hgqsjXhLIUCGFwgE3ffYDsyHIic2keS9Pn41p8roUqZqzuR0olgiy/1CetUCK/P73OBkrbSKOH7m
jSP8Laeb8FqEF5F/8ECoV4Pf6zWc261F2J7VR1N4D0+2Q+Xq2Ubz+Pdn9gUUqAKEzY0OYzhvwsV8
NucJBrJTqPZC7nXjyrSzkMyVCMpyd7Suv5Hufo4PY84Je7g40eqle9cK6gaB2yGK7vdZttl0HAp+
jK8SnaeAPIcLwVhan99hlbZRzQfCRhb9Av6vJlY2bvsvfdN3ug64Q9QIGV/1tgcCq/c0AufxEu+I
Sob9z/azVukD3IERnLcoKfrwUWQqHzW0Cyrju5/muS6UFJSGslLiFu+8cZdCZzjLmZc92jxCdJJg
hgDju8Sg4o+wBjoW07OPUDI8s/wIE6x1PcPSQBeu9IaxlBO/pI6bqyyb0mHOTABpNY4Lq7XSlveY
ao4aXqqsKizcZGATaOXmcettciZX6Mr0YIcUFf51FdTZqtIexmBI1Ff3c3PfrgOuAVKCJ6DiNmNR
fKxImBlRvBjzsTz/CYyzpmYYyrbO29Y6HlcIhlmq76Czc5IkYTviA3ZK+mrDg3aWSWcBocVch3SX
D6l4kTgj8+mQTpgNDyYohFf6+4IVZDQrpAzeXJexoe5UuDoAKmNKu9LH+K8fCU/f/8yKAM1OZsg4
S9k1lRVsDTEeF1KZNxnx+0FKLO5Z0Ipbpyq2zwybz9gO8X6d4xYEzFE2vkLAh8f+mrKLMoUJR0Ru
stV2n+dMQjvjTGGJ19sV65nasDV08h80F8IXTjfBNC0F2eCb2Ax2Q5LBBXqflms1Rixw8Qp4yeiv
WRObF0nzV0CxGT/z489nRoWtk6wfIko8T6BUNE4vVeuB1ZmjM7X3YHkBY+WXDW7vO6JHH4OT7QIj
/akzm2SpzCKd80cp6TECHRFYVPpmCga/C4wrdMP11TVc7NVkzzRGhWtTSODiSm4JKUvj7hm355vm
+O0mBHzw9fZBktsqFt0tNAzp3bvkYEDEj8zA51G+E75gdzOzCCFvy/hPAGwSHMT1w8OWSNUDK91Q
XZENtihOZRjQppeTGWWlnzk2gGy/Dr+G/dWFzesBkhIB26HrP9r68OKc48e6o2ftnyM7Dr3q6Pes
PNtxRvsbWNh6caKUr98XDxvx4kz6q0ZE9JhQgPkA8/IK7dX3LYCGD3BrhIIMa4l+vQk1w6KJxnQH
7gagJtnLOfS+mTH8ojrwkWJPCCXNs5bjJSbFQYIs+KB3HYc8F4+RcfsxZk5XwZEIF6p1UFcOQGmK
cvoPoPhfFdhchs0+B2wXmQtJ0BK04qTU9QpQhWp6V1Av973u2KV182Bqg973geAt/wMajrOAOfuM
JjG+GVqxD7ITB0NbFGg3PifFgWlbBDRmkRdkAYtK7jlHmW0TC9hn10E86wQjdAaJP+HQX988wvvt
ExRT4PQQQ0azmYx9IR0+SFQIcdjl4obiwyzKKioBdiYPq9VfVIeXzzEIR9Ga3GrMaE/+u2ncfZgM
FFN9PrLTmD2pQBL4aLQfDKjt9MzDAsXTZ7rrR/Nham8wDIDAPq57yj+c8WJXrb8otdX94imCDfjp
Me3vYTyq8lLBpjkvsEA9sLozesQOAda98uS+hEgvy8vbpvzeCqDLovsF9wqMkI4jal3b9kLe0K0f
VcfAsYu21RcRK+cXkhCrbRMoXB5yePT/awzUk5Bb+v2WPJZPWY1SGXTTjSgkuLpEOB163y1PlsHh
7RWGJ0PAYffOtCfT78Ed2I+IIJzZrNJmuHU1Xvpei1SoV/H+GYQq+/hmoG0iig==
`pragma protect end_protected
