// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
PAp270uJ8tcBLUcWk3EIy5C47eNiyUAzRH+FRnk+Nq3XcYm3qFtBhmYz8DnZR6azCJjfqCXInvVv
+kEtiylHihYFwhSzBe5A7+gES+15TLUppk/LEECakdUL2xsted7PPdCAuxLU7uAMugDMWGUQqKsl
acs3dztS9DMw4iY4UAXKeCrBeSNv24t9zHDJ4F56byncV7AL1LSolpSSgchH9Nd9hqY76DyffZbo
ib1SNfv3HRrovjsYoWRctv74WgVATT77zxkzJTLgbbNeVmVi5o1tKE86Nms5UD78inu0IPouR/vC
X4LWvpud7Hax745xwGt5zsD6bfNabdHdlvJ66A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22832)
DMewThsIj+Q7mwVrK/EEanikd+F7zyomBoZ1zjeh9ITUpxp2NnlWgn1XFvsIBejJgY0f/tA/NZMR
BFpUTr+Z1kKQKQXnCbbn1/fz3oz8Y5lHl5r1mEk/UCM6DNegThyRePTe9LULanSn5bkt68IzAAUW
FZ9OX57ayCMas1oUQwyqrwJrtdJ8/LNI1JnxrNv7/8eW4neeVttt3nlp5Ns9f9uqIWPDlJS8WpbA
xGPCqm+I/UxLpxmv5KGk3wawRwB66RakGfsCLtCp+kdJsBsZlkH+dzZC0W38M/IckismX8HSbBqa
LkYfA6DlWDwt+V1xiSoTHwGB3hQBtVeeGL1wBFBMymRpsl+Fj5wQRk8ymzJ931eU9cVpsbFOxYFE
aaxiXs/2foMmk7PtbBi4227ZlNCmN3el2vLb24lrWg0brOuvbxrw0wyVoUPmRrpFqmcGYXcSaqjj
RruO2bU42M/xqnREc/hDhZZOXlU7rbhYp9TI7SPEslmg9Oyarv0JsnmiGhB0SYyer4mf0dyakGOU
k0vxH2hrthkhH/rPxxaJY/Y6Z730orxE5WeXBv4o/x9UHUt86UmHPtJxcb9pnSf7jJL/rPqS60km
hpsw3YD6OI+iZtnZ7uInsJOYpwZSPjsXjyBU77K16LiGD/sA/wrktOhWyTojISKJGWfXudRbB/yw
nuTcMJsDFhx4P7E2svPibZoFYxbKiO4PsCZyj8kD3OaQkrYAKXYVg39eALz1bVkfrufcuZGL0Z1I
wmfoGsGmQ/THqHAWjbKmkFQfiYEFgwklnEMqvcuS4nDAWFjQ9dZBFdPJbaOGMpqAQLjgC47KOVKd
iHwpyq3Fpc8RYlAY+g+1vterB4dlS3UGM4eotCUDo2rTq2mX7/Uqo7SqbLqIaSq/vJt7srEW7sav
y8M7SfD4kO2jOTCOQZ5Z6mebXdyAHa4aSmThRVflc0xjBDEeQiHEG4N+rSAdD8Q/1KMgMrJkXFho
690TVf+GAWQQ0xwpWhj75WKZTbNrQMQPQA4a56fO8/FdTJeO51y1Ard9c8sEqsDFl9F1OKvc6m6H
Rv4jXQ7QSYqGptopwy8r6ZxDS+xSxC5LHBXGaD+uhiXYDFwCM5C/zh8le1/vtG3bS7u/t5HsTBvk
S8i2WN9oL9LTrbfMpF+da5LPXmscO6F7c2qwURhVT1wKwp+9Jelf7mkh14/s/2y6o/dGIl91zBqY
xoSHBMPK0YF4oOPZDpE9+dkp5BxjSRhEvRADtz/9He9f1b3AszaBe8LNLlHHazLn8ICeBWccOiRV
NjyhMRbx3/O4US2iBMXzVCi8ijyfuYR7KYzFMF0OmI34nTS9Sa7N5LKcP5744uWZ7RDBYkbwghMz
2HZ6DK/JqlKwRMxY4lSLc+K5SPDsczLNK2mCEotqLiIXdUCNy/xzyy42jaq0rttleCdqsjvCNa8O
j7ULTk2SP18NUPnzMfVEb5kklIJzT6JsWJ2rq6qLQxOlBU0Ar7uXH2roOJCwJDcS+Pfgn3CaCgF3
OKfF/+peKaC4k0Qj2wkoa9GcJlw0umHBff2zKL1WfLQuGYwdezwRajbzDcKI87yktis8RCl41hO/
NxsDpxVgMgCOEnNjct0ELLZPPcLC5r1m8ru1cNkl3q6d28W3et0qlNq2g/v70PgsewRhPRvk4GKA
Xdjux79dUUDV1Q7um4TSvhKopWwUbdDkJexy0yhVYiNWnWdBndtT1XRKaoPCY1i0fUb1S3gNpLpS
hOu8c4ktibpACJyfLYQza5wdpXiHVJlK2WU2uDbyDe769XcluMZ3ZcyJfbzM7+gsSzZz2VK8bJRu
wOOeUioLAH3bQHaP9NGdhkHUwJSJma5tsPfS0uCbt4lvYROpI2MVbsj2ZXE8V88Ti6+MsIiMBYA5
LnewwuF34zvtfylDneBEs8iNskt/Su1e+cksGpstfB+e+knw5J7FNGAStOqSIKSx5EfXPeTEqDz6
URFctUpGvVQZ3Qn6jOJuf4LSce1bGyCzoJKlgKKOZ+Dk/QPFp/zPxEBMvgFUqADB7GPAoQkblUTj
xzT/kwb4qEPB1mMEuNJMivOb6YoEOG2Tny8fhGON+wuMu4n2e7+LUiJXFE8Nj0rLN9LQmdASAdym
iZVJcsqTX/MZHiKl/QXXYb3jmQ8IAxUksAWMxGEDtunnMjM5bIkvlsJtbba/UD3yUapbW8zqNQNZ
ANnJrVWIKUrmwG/VwrmPMFwYNoiCYdO66sGcVyIfTQa0yAY9J08alfDPFk5U4TztjTHUwJINXrKB
ScejNtz9VCp+VkNwpgcY/QQkHqm79uxtG3cgFdOuNT2zy7jWDKTWQo0Gu/ufn4dMsqhqplps/P6Z
asEVi4/Nly9OLj/jIxtkXbPjBmMnr4Nw5qrcIRm12ceMzrN0lhaur1sUX2OwuRACJGFNh/2dweCx
dfy3weAMmZt/+vFadsLym2c43mx4shH/lbWLZs8KmwIuRRXh1jVWLA7y5rdxx5bJMiGBCBfLFhKq
CthoCinOw7LuFDWFDx+Ub+Z7hv3JyWBmyyLpSOOLYXpYNPFVOgw/+sjbaBa1pjjeNzZkWD9kXR+z
1a7IsycC7xkqicRmxnU5S4aGaQ6UX46e9TxWeBArnAKz+1veSqNDavxdnFUbJ8x4cRpRk9rczIYE
lk2yqoy8B8e1uCWElkZbiFTcwFNC6PGNXSfuS4BUG3M8KeoFSsvZMg43HE4OdN7n+VtjtNO6ONS7
7Aly5aPPTPFIO7HH0NiKUbL/iJRXOyvR8QYSI0e41RabodQinSZUwmf8WngA/1/kSSk+hRgmlQkZ
rsa50LLW2HM6GcV7BtDfEUkqBNUBeM7gymIE8yxHEq7+k6J4gDVDBe2+9N9ng6cdAXFJzCkcudcZ
nmhJinXSVB1IyEwXWXOzwRsWFzPibMLPTNJ2NoMrMTEOGmdIdHSIoKYkxc1HYNgcHtnisDp8Pyc1
+dtv/JnlyBPBt53pSs79BE59ZWirDE/XQgYcOobl1bghn7T80Roy03ADkCyhDPcv48unhKGbLdD4
JLnoP+DZ156LjYEl2q2/U/kpjJjyDeGs7whltP4/yd0k92L/+x84z4nXOIhtiboH9D+COcOYjRG1
tZgrmmDPRro7tZovbQzCnAA8SzFCBP4BuJmcT3puLrsceZSW5FREcOVYt3QQNc7lr5vXl8PDV0Ok
QeeiWnatE4TfgEf0JuJzEcoJoYbwZuCSLV2f97DFI6OABISM9uLayoPYracsPn8nbd3l+LzwwFd+
Mhk91R5rQ22Hhf8Xu+IOk+y4Oks4WEmosycM1xCEC4cjf9P0xMDI+9WWKKaKBqBzSTzFQcMOZAvJ
kat8MUrgqpzUVGBCJrTMCONuG3fRO7tg1B4OLIbP1nAPyU/Dm9739hmtgKR9n4dfdA4MhFZweN92
Yy3A6J/DWDd9zjfKb6zgvuXcvVOJOQVmi0vpAaMALZJBLNAWTX2GXvH0iajQNHCfsrkhpyc4O4Db
oqYa3pXhwTpeSch9M0r2+LbmpmkmmBHJDHkUwAd74fada8ag76v/WMdCIVUAYRAsOwDS5TnIP9Tq
KM+AMH2WXxA6hvE1aDfVeS4ArGJjkdm0UglwjCYhzewLLCBLmQ3XsrdGcmsUgkmH311gZ0DzdO7Y
mpKOMltBugFGYQyh44VrppZhHM9IAN1xuPv4Z5P2sIUFK/LJS7QmpZbZUROcOFbsrPJp9E3gqshK
dhrFhdHo4R+abk3BgkR8impDhwAoP8RazFSYPNNnSkgk2kshgdf9HBTUKJczGyPpNZPH9XDaFaG9
9f6Ug2OX2HYxJKZsilbEIwWtx9flNBV6ITMA8rB1yqLtZLT7Zce9GlNmh+ArbW0L7euOPvoatmZb
jFf0glJzCBBReFKH91/Rf/4LyGzAj2aC62naOA0gf0gl75YKfRbkOlVW7QyLBFv5jDhx42Xu4AwF
2cUjx+Y0D+A8lnWNdrZn8ifrndMBnDaHSxZ/lvUnC4o5uM5SAcgRzM0ipkwNXcViVlhXSDhbI3uJ
ETCnmzVnHwTCXO7NyMLEOn/jqFS9z7hxUNy+wXl8quzSMi7Imu3cuSwevqftMDvCkkmQ7V8l5YBM
YwECpPd2Lg6/TsJd7lQNC1Le4+lDYWoTm/7C1ZhYsIs5LLJenXRrvDZO+jdHPi6AW7I8UjZojr/w
xmI/JjbxxyE+tTQmtT+qgtHbzb62F3QNdJlAab9vR54Rai+p+6UlRrSX42F9o/r1Z2Uidxddy8m8
KAfqdioBmE/nlfiEzdALSQsPtmiOKQ330yjO+kjhbsUL/l5OY5AmaoAq1LHCfzsaOTzlrF36G/xk
PuvICq76IIj6+r8ajcoQ7I3AT8ya+D2bBTzcLQEfhuieAUCQ93zPuxZZcKl9Jg/1rLyuqtcYBrAh
vR2f1ncgyO00FikKPTDF45t8VhdrI9wtwnR0GJHwKY6geTGFRNg63Xpoel2oqZr4bSRkrBDsJ1VL
/gwiOQrO9KH8N0RcpYWcufv+J55yUrIeLAWZz5ZlNzcUHEPdcEfZ8BuKuqTNzm9ycFV/vL0ScwzW
Pp9XNzNpH2t7i9dMwlZ5KZw3vohgHYAZ/iplcc5uTE+Wlr+xqrddYVL3JI6BaaDZLcBudgiBY6TQ
qV+hpc8RvUkACqbVyD7vvAi1gyrU2Cx+t1BLUxxJ8rJ5cgebHpo8OGmfWS/ESQwF1QsWM67knyL5
p0VOSOKso64jZbEYl6+mnOHI5momK4uQY4DtwhvkdD+rvINdDY9uQT7nodnCxuriEfpoZnE+gCeE
zezaSP/OsoNZbjc2VWXcDgsaz5RW4ZKFBrVKdAyVtc44eOQW+WSKdSGwXZD7Ev8vIQheqRo3+JN6
sOPmS2o8dSk5D03ExQERRlKdA7yb+Cr7Om2XuNEffsOXlcSd0iK1z9KfLTZniazcHMeSYWVFuwBv
vMQAGovcQ6j87su+J3oB81dQjG2z5CUxjMgsk3EtK25tc8IfE3r14+B3IfMMI3aINxSOXYa5gEKC
D5dG+0tFs5UhrA1kPcRG1kJIQOVeyVeakKE2pPEFo61c+WOdKsXFY2kRGFAZD4u4elOJdDf9+xen
MvMo4f/mEFet5mPx0wvUsfUCL++sh8nwd7Sjmdr0KwESV1D8+xRj9PmEWd7Mkp9kD3mUgxRlV1mL
shDbpSeV2OFMHt55uttJl4q81bVrobvXvVMldh5P4E8J3ePDZRxNwulFEiTrwg6jb7gUHNnuQUfe
6/mgCdGNkCOKTcTyxg8Pl40PALWHPD2aKT+acHtFeyjLHlgDbQg9QXlnBcgTQe4P0dCOhJGAIWEi
JoDtaTWkZDP9sES9DJstARxfoBYgVgnFuCK7KSUr2QxnLtnXjMG9983ZfrcYFbhD0Y6/6n/Eko1D
U7b2YHyCg8dmSZ/igILrZqEc/BFY7K6OdJE1fcuSe/jRpyU4q1egNJvZBRPbRoS/2gGj36HViIPs
wy7UCSlqHceHyZB/SKC3nL+P119jOxRkGhiwiWNU45cg/trk6T6G21DCfeUvQCpS7OjocEFrlpj3
E1A7ZVM14/EX3rZ8+lj7bcu67Hd9ayei8oTw9IyVjbFBEJ1J0cmpgsZ4nY3FHDyG7f9ewLAS/QWH
HkkfwGEXe+bYnP8FxBeitgJSeI4RoXeQ1Y+4MbEaKYpngA7hMRHQ+n/OdaRfh44OUaFEW5AbP0T0
FVIa527vVtXESXz3gVOLSu42hVFoeIs/OxqDgUl42Fm24lPmSxyIualuFuNfqD4Jkf598+S+pmHo
QJoY2C1/8WcYzqXPa+e2mUdeJ1Ni2xdW9WDHyKldE0SyxFw5hpSH3VJbnhbfVQRkB6l8NQpGQ/4F
LLHTIsQpc7lRnT7Aiodaf9w2Oee4tJorGthjY6Z5S3NRNS+UHd/MbXUUQV/Me7ZB10UwmK8CEY0a
tpLGO2OVsZWPh2coqtGHwQHYlVlANLafFp3p8hGX08D7bKEOAPr2WO/gGuhdn1v1N88R6jFPifO4
Kgo0RPabpjRK1b7hwp7uMXg++VPWoYELP0Plku0lKjMBRUa7S/c/iLz9Iquzki+7U00rmp7DG2Od
pgmeTanzblzLv7nn0hqjIEpCZnh5TGoREdLnnJLOROvAdTY70ExjTEdGm7chTYn/fLe+IddB+Dc+
gsZIVtrUOcCHC5sbdMBaCSAVWkyTtmpiI7CA1ziKEROIt9aXGw+H6ms+rOOosOxHdpNREyoGAV2i
X6rrPOa0AdRU4anHXSaRiuEdq08/7yMybkLXdD6D3Frhnt+MsxjOXhbrdhNSspesNpz9RUfSQEGz
9Qb/4mQH1jT/QSF0PLs3UXr08YKg+aqa0F5lkCVe0NNeXbGHlsdZoAIgOuOgjeh6ZauOH0NPXSGQ
S3o7ghduYX/LP2xQ5jB9d1FF29g5MuMwt0MAZvdlnK+wtvMqguIH2lfq0Yj34UQUkRpI+ibuaKDh
WdK3Qtrk4oMz/RLdgmknGaoCjnEUbRl/2KozlZEkRjJoqOCpbqJPg6zbKq9gb0CE3yLYkoAATar2
VnBltBkjNaEAKUq6hIE827z91yhXar0lmMTDoyy28jyysWysY/FMwjn2+dQoJIRCTYKpvkfh6Hr1
h8PylFelsI9yjNwGxHHnIRK9J4p3fFLCXsgxHhgBP9iW0xk7xnNf2r+9Rcq6lFY/zAasu4P0iRYj
AK7kg7DiJ1zW85hbSmYREXtkYvow0x00XJye+43UKO2yq29JNHKoMjxxHPxUhGaDYfD48Q9A8alY
lL40dg7ZC20sHM9FvxELutWE6qf+tsgacBfDRcwoCs/MkeZ9XCxjW8i4AUfJoZABBF/wUFCWx+p4
BzMb2uwxDSMWAXXrTerPkV+AZ3vufkLQXNx17JFkyPPZUHl0hCJjQqieUej2HROau5esrrm5W6nX
KFW2bLQyJbb1U3YTPUT9inVAyVzAJw1GC/5wdTHfyb1a2s3NSubSajKPHYZ75MxgVjFA6QuO5k2F
3NrU4Dz8+xwyY6mNTrxdfaSi+9njqkMnpS+ZqMAgYRMV449yYwO4zkGms0E43RS4ekJFAu5+lKY+
e199VdX57F3PlxvRjxlJLqEgcIRDjjpl7lbbK1+IE8ja/8LIO+5ZQNgJHpdm5q6xoRr2LzvLHrvB
LuMhnXRM3gw/wohoD0p7htGoUy5phLa//EeTuxU4LWoCs5Jc1K4yhK7o/RuNdnoHBnwM9RhBdZvG
mkMKR0NmP3p4h5y5jNicdtSlW74R0EZbc9JzafHcS2XdbSQzkl6PJnP5YxogNaaxnrKCN1G3RvTq
McsHudktLpYR6bdH4vfpX7d0e4E1Jpn9IksZ5v3jlFNy20m8xXrHHCnEotA0rBdWUFLxb13H0WKv
FZbTQH0WeiV4rhHTEcw3pdQB1CmlLVUh4yNkOz9jxrX8Wwf8sQmBirJyDNt3zxYBeX8J0bSmphV1
AbvdU9pFsUVbNRTQnt2FVeu/maBtlcxhfS/beanQUynPbU9ZYVBQOJ8HQHgQkLjVRkrKBnmTVT3Z
0ZAhetsEhGcEnROeun9ImJZUSbBJwnLrOZem15jkeiKXJK3su7/5aNY6RZrbNkM5zNfr/fJSf2G8
1Zh9q3U9AyuHo77gEkJkZFJu9tg3QxZYaHJA5QtxwCDn2X6qQuZhbPHXuN4PPNmndQz0QR/SxNlz
Hux7jFTs34LMNnTWlVN/EwbYFNjp0eccZt0H14vQWaDmek2T/FcIQdnbSlN8/eDnkhojJC1rPwH5
+XikB0zcPCCii9Lbw+/UEdqtA8iGpGnzUr99ppXffw/ZjL5HiaPdVW/P5HMBkJrDu6NuwvM+NRVB
ziTDTolCuvmDBpw6HjthiUrGDQQVTVWP+1Isz+ErzXY5g2YZZx13VW2htJhQn4ZokPc/jtREw/NF
/MqPETZ6DfOrBqoTrRRmd9Z6ly1u+p0sd4uDAjx/3SsFtQ4zl61K7wPnCrBJZ0MUA259EOddOiWc
T7lJ5cBBW/sGWoIP9syUkCXWtgQJStTR7ZFio1y7AZGMIZefkpaPCMUwA01nvJG/cIX9aBFcisYL
zq7J46r6rUcT2wZUg/GfDg7DlemXzZukOSSnWC2TedrjdlkJQ5a5GXmfAAdh8WzAfVYyyrR0yfVf
gfiZ8xRxwz1gM7tn3OkZZYDw0R1P7h50uJ2PGJlVVkDwgAwAf9aZv96y+AkPrZgXKJzgLTd8FUhH
9oxwMvlD5YmmbQytiKsn2xV5ahz/WL9Dhap+NrI8YNamPFdgHnxiS4IYXGHTaXW3EEsvqzlrMLW6
c0JXzHLas8ycXwm63XzpM2CaHIYyuDqXoqaOhAUDCO+j2NfkVMN3wDEW5TsEg+kK/3yoaguuoyTs
rBha5BCASheAPcAA8C0ojbDDIFsRWFe5ya+PyxD/+qcUbteEIZ0kn1SE/pzvGvaqVhsAz3u/kg2o
s5ZOoDgmLmiiixI/Hw0ctU/ZhFV5L05BQtndLWIfARCXaQO78bIkaghdmOS9jRPzp5Kg2u6yBj/k
Cqmai0o2mtqKRTgcPo26n3BcaZFkVzORcwI0p+Rf+2hHRXank4Lf7FaQa5BC6o9fTcu1qNzWcYvk
W7VRlOXJ28TWWyz9rwwHMGA9MppGDhbEzqkOYtkOnSy12bsr1HfXofcGxSJhzUwyioXZj2mckSl2
z9rSwjRRYQhZ9s0Dng4CBoE8GqxiBvCRYskGhoNTdsjtVUNZCr85m/MVj+FXYSB8YMYZp4OAnLRC
ZPAYz/cg8wcxHAVDk3CHWH4S+MOq5inODDLVfwPyX6U19LOJ03od5j4QAlPLfJQycLcmCpkMkLcM
aKc0fGeREV/Ikr0hLQcTg8LboTMCYRZYWvOoNIjmYPsYU6I97Uww57AFfR/ZxJY3BR4mkHufmXFi
C6A5KAlEEBrjqhCWziAyDq6SyTpvosENoNSnlxWMJmD0t1PZZf9sPSgaBiU5qKAGl4S/+80XAQdw
c9PSrcEgNojRYbjP7/2p4iR2MvLqbCCRIP7OpWuZuiXRuiUQzxvJK2tCLoC5NLDw8G2I9ybpgkty
5mlSvGGy3DjmH+22fgZh+JVwJeyD1WugnvzErrIFxIf9plp7XNowKg/0Btj3RffpdO3Iv34iddPM
W4MZ8KXBVuR2Y1yrubS7Vfae9fp/LIOoo4f4Wkx7Yka7i28SwJaZNBBiUfTz8vAV0klc9Ejn1u9e
z9WNdlnbr7sqq0lst5IlJWp/N2VD54HYf2TUeHIC0ZdmM0JXVbMuIJw9iCuo/NDW6M405Fzqajdo
kTKtBgLgfa2iFSmZ+wHer9KZWi5T04qZEECHDw+JNxA4x4+cqeyM7shClijazLjpPgN0lAnDVJEP
VY4uwkgF7AOKlfcKxeVDWD2swMledd69BC41JTaF2DanXP9IYaoUAi2F1wZQp+/VMVRfW+imKNCQ
o2LygR8kD9ds+2OOXITWdQR34QSwwDod3bcu04KsjFiGwUBjbRfgR3DeKeGM1Tjo16h73JfPRNr6
yFHcrG7wPLxiAcgkouHA2LKd/upf3vQjmoQtTz8foeo1VO70f40GGt2AlI9u32Rv4FXMP3MbTANN
38SYeRmHNBVKdJk7jPXQXmJUERHbKJbgdRlJZm1W1zY1rwIo9vaOGQ73E51nkq5f1pG9YLGb17OW
5QcNYK3fmIomDHEDUuj5wtFfIBFTZSplrQV+Q097yBhYQiN/HrWTMlq1MpDH6kjDvd/+cIm7oci4
U0QkyZNv+1DpQN6ljYMKkvTvoihVnmqTIPP+l4xZVHk+mvRHBD+En+ih2iT6ERA3JC4DmhuAoRsn
RzFt+z2lHbZmMcBJSceT8OQECCMzuwR28c7yNb9JxkPWrNDnBZZMyOeLRSmmKuUtvwKRIK+wByka
o/L0seGDDYzvAZWg1W+d80EYplaOQLWgcy1THM1CfkL0pP1/otyX3Ld3L8viqSukTn4c6ml+5lNZ
R7jquNw4hR4smIuxUlpOFFydp+DVn2Z5os7O4Huxu3YFlR5g4v8Cdk3wAEy6wZQHXrBA0G2Xzj2p
JWDee04w2QpGp6fhOOuNIvVM2PFeGqMAghe8peRlxGNzg4jTFSEOE94TI2921nw6vt1UmyG7LbmE
OVdTCshGXqtdIM7WBToWu9O19uDUbZr64T/lhjcoxZ8p0cAy9h/8H7/o33IaTImjPi6PaJ0ej6LJ
LJLXS0DOrbCLmVCv+5e/I+xX9VOEBR4oIFxhAY/WrgwOaY/QWqw3M5Z6Bml3ul3va4gQVP0z6Myi
/xt8nvkmIQw1N88AuCEtkcKWlghYARe2KK8dhtaGJAin+xlwFiv99CbmOfs4scKm4edJwoCZoZSv
yJXK+JftB/a8niDOp6+IwrrOceCB4wuEIRnp50wJ51onD1+CXa+6K9btNh6C9PmpfQ6YW7dStOfl
b/ej59LcnI84N8evCN7efq98+j17/UEq1nWPQDZcWxvru2pxP/6l45URvL1yKKYhkgPdjSzppqgd
NX54JYOOD6U+woCu+NHaZjFC88rzk+pmt5w3nObaKk3pxtb4M7ZCLboLwBzm6R/Ck7yd6XGc19CL
YG7ySynkcgut9OnJ+hj07uCoCFgAc3QloLpFUpIjPYfM6HcYDGX2EHbxXc3Jqrgxb3C7TGZtqnYy
fh5lExVzYGWWD80qFQD7F9mOxXC54K5LAYeQrGUsyaYo6YDFZsVun05dIjh5ttIltFbK7eCkDvWB
6SpgeQtQUqZJX/aM/7aP2on3c0/EKH0xPHkMiVETEMDQLSZt1rPtgfqysH6vPYq3W9sOCtNNCrmu
bcMBXcpRLXxWoqYr//v961xxD9c3480WLRgIwPnaPeWOk0YntoJy2+dm02KLDrtCy4gT4XPZP8jl
KdtNIulga19NvWKSZQdQQkWQO0L1uCY3VE2bNk3yzhKBzdnTlc2tsEa+jfYW1gHab13/N11jiIRz
r0EPPQoDThX7+JSn7PJFfJ+RuDfPgi29FZHdHdiP0oHMdlTDfCWbrLZgwqgjQ+XKF9uHU97WcJoO
beBo+4YzV7gI3K8zs+FrFHrqKKZhOdpCurxtLwqe4y451d1CxPrg+qEPZ5j5DIB6lOV56C0vAbdt
X0Q0itSxqeLEsZnmNq2dh2bzptQhfqlyD++DithgJpGEEj+Ein8MgotFdNl8gxO0iwGmsbEdyAKb
btnhn0RCTJ1xjk1ucd98fHhZSBEeWH3EDkd+i9r+XpcGttNTRdMW5pkVyUAEyflGFs0Zi4aPpjBT
QWCAhuZJUcAEQvBh56fuQKa48vrB+MeMzVoVBjGVVoniFfXu8kKfeyvSDQcyOMXs1ttdt9F614MS
ZzsauGv7w7tKBd5YMkSR6RSZgQcop7j21+9SvbJlDlAkZULc54yiD5ioeyZACoig+md4t5oBkATB
k5Y9HIRN0ELdjyW6NIaT2gj17dtSeNz9ITxtZjDC5DL69D7wKf4bB9vw1c0xWAwMtpjTy/lFFkEW
lPynrnrj+jwBrFlADFu8vn1K52/sXH2mUwo2L0AHwTXw+kdThzrQz3MEzSAi7wDjWEJv4Vu7umvy
AYz7lvLLmVODt/FsJ79lAlACD3KWav/uutoh6AS4cU/h4UBP0TgCBQp7oBKqI5sLs4m9+yLUSd9g
UhbSIDtiBXJAdNwWF/Irl3HnVYL/oUIc/RIwrAmVJRATcXGyatMfg+I9ACR0dSV8pf6O7GZd5n7L
jfJOsxcjupFmlnP8+a8xpmTaN9vp7ZOsMNeUwEWQNCR+PxnG+kJsosQojFnzssw5/6HqVEKB+tIn
guGSSMS8PYToG5Mr1AXUNNOlAS4nbrXG8DZLj7nZEIv0GbbN+qoKJjirFevDRyD1sBZZrp8PbQoY
C8Bxtv3aBzdRweMpASUn119TiL5NgyvFfDI3ivrVaiWP/ZrJMt/ljdFSHnwzf14aXENHPwl2DP+5
AT1ymtEOQMDFEHHyxBe+PlQQncWza0bnh18Y9oKAkp2vpo7A+n4giBn031IMCUENiBXTdKTfIbSf
sCjo7KVDrK7ry0sZs437n1FrKwJLLseu9E1Rg7N0teqCzcFAUd/NTdqOqRS5oBb5DMcdIX2+E3j6
KSzPdqo05pkR3CmuBv7LeFh92lk+Z3KM+7+hWOjPcSVyj7OUyblzr2y9UsVOe1WN8qknkNyvcqK6
snYiUOing0IlRM6RCNweEVbk0JIyOLG8xsadee/usK1oMyTV8FlS5JwzAcEsx9UChjFax9Vfc+kG
1nG9NDOaSiCfXHAFpNHQMplLFA00u2B5vQzt/nmo+/SVO18LsCzJWYIzjPQs/DyoUJ3Y+9TcJLc0
YeRDIF++f4TJokx4ZPq+M0HXGq44029/KI6GWyTtO8qKRJGDPyd2LZyRLyMomal9xelCCPcnvd/M
TgR9HoNRxZ/HfU02mSHAw2D7jsK6dGu6DxFUcZ/nMkFdUsrO+70KL3isMbuJgObvFbl2Qt6eMTah
Uq2ILJlFtOCWrCVNfoi2CM+w14qCpuuMZ+lqiy8bvg6fIeIF1innv3bVPEt8ObyIuKlHAgW+4fEO
LVuJoKoh1YibTaG8UhH8SSMlW4uT+TTu8ZDXFazhFzvQhMblpuvPDHoVyt3v4mxFEUVvcN3EW0IW
buC5NNMswAO3ij2kyfPpRZqNgaMT7ouA4mKiL8KJ9PflgpZJbOb9nl2ayJLtQozPUSiZcLbTDFjZ
BDU2UnctCv+l4IBcaWSCgs9rxC1tBTjuVH/xhfSEq4jOojkhSNni9aCEVpPspUEfmOUsZdKymPsd
49IiKRdWEdNhp5afisRIVWyVskcm5kg/TTKIMw7MtdlIf5k62WEzH2mjA2k5wq/WD3n9cXDHz5cs
frnlljC2/T0jjMhpVnh0hcQkWgVDCKJJLkIpwRlbjrW9iKFGgrarLxw/eZC+w0V1CHEHKXET7EgR
KON0nq5TOTyW6AemnDVUFJgKQzb1x9aNsFnr0DeLvZiB4fQPcx01aZlrRhoZkfqQiW/jv4HicxwO
dC0TUpmYtc+EB3drWqboPh0xmT0hE1ORsno74wFJYIUgjBpNgm2WAl84cNXylPqAXD93CDN+R5zh
1ae8O1HNsAYCCHayMIEAIgHG4INDYAmAT1A2pVzZB3UAxWomrXgOQY8Q7Y0y74ByeOnpXPHpnCeb
ChW75xS5ErnIW991xLSyeKX+obA4YwYn/xuOSfls8tXr0q9aC9Jc/eCqoKTt+j7d/T/fB0OCXuhT
rf33lKBRguaF2aP2alkP6JiTovsJjD8IieifCzAO3U0QHoo6Toxw0sifK8LxzwxqNExGBB/H7P91
tCuNqRSewzDwQy5gKQGYf9xHxly+nJdOnPTxFE03qxvM2J6ipjufSAk3bjRczldHljYiQWYKGj8f
Ax+aKafCmaFzZGhbQGUb0DSIDLDBTbOfBUmMsVEbKxLr5yanA6sGL+7va7L9+SH+DTCT41xpoLC/
+YM8l73ANikPXW20LWZEaan6oiNqRBdW6pxvM5Axl1xZqbA3cMC5okk7gC7dfTsZS/ezfIy11D1O
HzTtmNSVzzy5wLKuU5oii5yEUc8rIfns5EMSdvTTZwgF7t9d3xqqzmnDO0XaOOYyaAOGZzwAYXar
ZeRPcI9Sb6+y2HKeGVV7VV46QV8SwM6Pzt7E3GzRmPhyTGPGlc3I263rve60NfllZmyC2GKYCJev
x17iAy/sO6aXhCK3fp0IpW4ePdJiPuvZqTQEOls549zMvhwdJxdKtjnmz3gzYv8SEpz6+ZXBDA1k
JU6WPd5OApvA/WttsJYM7neDVzcqQy0LVXh4XdcGVdj2LrVr7NBEGzeT7v5hrS37/FH0L0nf0CIn
xVF0n6wPFdiyarpJHQ2G0DAOfLsRO8sK5w/09wvbOnflQJ/7FvkClurutRlB1z0TTSnDvx/sZnmt
VhzSFtWRWGOY8sglcUEta08+r9mJl7Icnv6plCSdyG15e3ZQs6mou/fmdwyFNzqeJOfa3xdUVGMj
mzTI9sA0d0qMN0KTTZ0edKtdZoXvx0FBpg/L7QjKhGIOVZ26bLl8SdTWMijEP6gr0XEGDbaZMDNK
m6XTuShq1X34gkH6Wx7BZLufwsVX4H/1J18BMvO5EBsTOj+aP5QIos66cTuBJzkPVqjpRy88aqbY
ihTQRwwX5iKou9ar5DeHhT5unkd8Vc7TIHml+KqxxhCbp4sHWQE4ZnMZBHHUiI3ll3Ju6Hb7HJ4N
P68Nv1tk5O5Uh0Pxji43MWkFDLCxAKzd5THljxsK3rJ5g6eeLQHSFUsd8A5MMbHoxn2KSMZsl73P
ywH66Lxw2TvrUB29KM9HU/nkbF2R2WNG/TaRgyboUE29pwoej71Pw2C6OXo34ZufF3ZaBSP08Gcp
x4VP0graIu/R/5yW6EGR8rn1HfY9AZd6uqUGE1yUEh4/xe+h6I/A8Q89IYiLfHZ1PWAA28tqjuxm
CKUZRq8nxA24wca/rckUQX4Fcvr1ixauPq/O2C0wDYVszn9LARpQlQNTwKGHmvuDf8hfVj9ZJfnw
k1VGLAajeIJHx+upQCrKL48DscYFY3JHSJy3b+aCug8U/5FsJoyBEOf93SH968YxaiOLB32dPJBi
bOWW1wpin+/2WLksKEcgN1i61iK4jaiLZqvqdj/eXETkff75TMxzwjpPCIIbqO4wsK1jPxKP7dNh
IJfiGc/dnfxQMluPYqGzQsQq41FAG6EkJEttW3T7XU78S+N/ePIlySNEtGcwRLaeESZOdNEEP4ye
dlaguIPyigm/HWUgZo8FoV6E36Srlc6oLuh1+d8AG2yV/Af/LZV6KBQOFiqfjYmYZdHB7O6kSzWc
S+hg4skEC0GLRD+ZThKfKT4x1qxi//2Ngh/uAEAfcrwKKlBUYl6p7yqdMW9THUp+6O+40NN3mIDH
Bp5jEk/ieic8/svma1ZXY/ipfIyIpMjfbvUG6sXYUyl6PDFBEibZkwm0Dbeo1ICW0Mwhwe4KEjlD
OFK7F1fJHVFOyW9U/O7DVV7RGuAsKOf8LYozQgPEIGOB+tGkvdHe4Ag01zPsBzrl47cVjvNrcAgH
d4xrDUl5VC3wuiSpH3B0/QAfuAEOwZ/AcmBXab0/wZAdfmDS4OTurLgANJR4FsiJOLftAapRVxIP
IUzqIBBbblpylrw+KIb6w0Fe8iESghcXHPM6muOM6uBuHccX4ms5HybXI7BTpvq6dnmPNwcMiJAa
dX76lVJOOfL40x7ev9xspcDPdiwbj+1lAv+fmBhUnJSu6mAZXfC7SGMA679BVRZ2h/bH/8x31dfQ
bEHuyWKOSJSpWsiILIdKYUwDLwSAeK+ipDrsZR1XbedGyP6jbQfDg72oIkTgaBJlgGJbsUtWG9eq
XP3oLOWNLTw6VtQAe0MiYqfP7mrQ5swjmritnM3MLThJXXhSoRuZex8pOLmPVI2cRSYcDPJqyy1p
oiQKf0E0rS/mLB8kaoBLQ8TtkaamERjY0pDUybDe4qt2yB8Ox6QC4tWUSSkb+fp5lg44jwDaVnIp
vlK2pL4qJvlL9PkI2c+ulToij5HLh01ZD8JsSNxhkUUurtvH9aofOypmf0r+NA0IXTndE43DGYY1
u2aGfNvOJR8fvQumxswzckyEzHHcshmflBca4fb9c+9WjWgYyaT1tKIT4P0o8jyCyeufCLYTPxEG
EqFleMJnsTY7Rbnyrl7g0+JpksV1XzQ4XKyDgcYPdiBebv1KBrBNki/zpGjNy159EnG3Bx8kkXq8
m37iZgr1LYsC2MfVHLdIbcmiETcZ4JK4WNUa8pur2ukpLchwUNbcO0tN6qnge7J/HnNAU11AidLW
CAVIjCEP7gSS9q2GxmHvTyjn0qgjSJ3E0k4fEsU21FhXuyADNxHAqFCPgqzqMWXfX+oMveOG/M4o
uj0vHMIeQfdikQR76ZOe3/zAPbGwO5E4HGzVpP2300O1BO7ia8oaY68n0pO5XMHVpvM+EMxoJID2
3/CiUR8ODyyJq+RzJzg/qYZnDF5L4ENGsVnYLf7Bg3Y/IiPLsISrnu1xTfBHxUUOwkpXGzGv7y2W
9d7H8YfOLRzXNMgB1i5g6KqFFzO5ckdVK3/jB7hfoWrD46OuLvsTHBTA/Ta9BjQ38jEJEe8ofBlk
JPWMF/+Pb++Qto4/gTCPcjMLKOUr6vRqryocZu8vp25TE7p8EDf137w9Fx1ktd+fEi9BZ56WTH1+
rY5tt/aKRO8SL7LTDpvUGQtoIiQw4ntWYZXPE/EP1oz+830SuUAkVZ+9WXPATtf0KVssEP0f+jY/
+8mucnkdP4ZShYfue32c7le0HGyDCn3QsA03KDq6F5OQFx6bag2tqYUNL4PRTOGQTT2f/cNnjPUK
XXRVJ3tE1fsOi9pdnW6OLyfdBNIxA8dKl0gO5xWuEeY/4aVo7E+3piewt8j2iUf6L8DssjFkOWco
ohL76FmTNxKNOpa2n6eIyt2DIAt9bhaK9azCMVv44mQszW9braG7RAOhm/NWWrqR2TOD15UfpyFD
r7qW3vzROeGMIio9hZaMHP7jfiqIIcrvMlFEcwm+WZUEny5lFi+L0l2ppHspTzHPW94erNQ7uaXh
38GM9dKVY24OAZqYkYBjMyVNeRHczoTLh8Y/ehaklanaH3HiaM47QmN8VjNWmJLUlpZO1eO5XJ7d
xBCyLARgBvtb7c6qybk8rqBcIuGNxHmRpOQgIHFyNDcMcEkhRxq0txvo1XdubfODIdXY18dGrJ7F
7qtMbZGwPA40Uk6O+uDmRTQmRq6wRGnWXAJ08JCSUJuoBbxW+TTkq4q7AjvonADPtPFvG82go2uU
KRvcvpzUWWYtMXcl6iQD0rN38KyZyRnySqYqtsX+iz2F/RFw24ltWw4dCv9kFbxLAA3ib2xnfFr1
XzWL0Hq8VLMDYn5iodoKuEpVFI8kK0wooFSwnKlhLLAS7GkO9b+7SiuhXrPBWftrMFjhN1bEy6vV
Hdr/4OMnx/A89ZJ5JW6CD12nGHQcWmV6QS9NAlZk0XAHypRfyk9oV2QDBOXLN/OCAJ3aKnpnolo/
lwGTliyU+Nx1mJcd/ooCjpEHjz3jegM9d66qKwcHv/aNDsle8zxtfGV7fTRBdLX9eO3x1wnGznC0
QOkQYQuuz3/KzombwIo27WAH3lOUosdQioD5lPm14FEhxxBDJ+FYfAT28JuGZ0iRLMJvTvkYsHEr
ftPj1+iwPSgFuFs/qDS3iTgPpvjOAqRKR8T5NJZR0f+5sTKyLmS6q45Qo6ATcao2KERZqj1DLWxF
m8bHOJOgLE0klxm97ujmpOfbxWu3hbuBls7EGSeHqkg/d6m3D2P9zR/yv2MZe3PdMIUa5QCI6raZ
UH1sJYGQ1mkYjiVe6hqcEXBRglhxVF8NYd+u4vhPaMtfLSZhKEyjBzYOfBWsMMhUyP12l4SHI/Sd
wouQEP3r5+vyBufIx/0KFYouOR2SDSuG/0m0fz8PLDOPB0hal9Z6uZqF6wmJTVY8RTBMKmwLdlYE
Vaz5ATtQaGcg2pYydey0b7lcvmRYUrKATI9TbZjZbzOs1K+I9RGWCt0jXhx8l6q+UD66rBwSNWRl
AyoE3VHHGQiyQsVkYZmixWKXqsk408az4X0oaRXktVR5FVL2vnnd0x7PJxhw5JTXDepRfCcKH/iF
EJ3vWriCKNId7ixAPpLLbM5GMQTqyoTOameVsJcj3zoFhHB6urf6K69zcJ0/NZPsyNF5G0ZXVmZW
9IvBM6ZXny6n0pM8GL/SvOz7SeZUytEzwSqXKHl1OEbyBbUC2RcQR9At6wKGMkKu32sU0MhzmCIR
GxhJBhMWeGMBHFQlZY/DR8uYbX83mrge7RpV7f+MNpaqdhGXcLb3WEY75oNFGtVGHRFs9vcZr8vx
hEPAZgJtaOE9CDLd2tKYoISYPmDif5/xiUh9bMjXhTpF5drtJwtQL/PQkICq1dq7tyMmcXzy5mTI
oHCf3d/Pne3ffEcFaVRLnKOxAzp6pUb3ERwMMrehGWYYe+YVLkD6ooQ+b++dKgMsPpJV6oS8Z7aN
j/8D4j7GZ2DsmFO74dmQBnU+5tXrnDGj55RbsayPk3eTJxBntILUATlNLyM4tRdbutQ+6Kf9TQbD
uqclldI1ayzSdb8vUVGFuO+ZKrqbx2CuaCARw30cUbyy9ftDK1r10fVsXiyWC3WA41/R4Vvh5r9R
eT7NrRIBjduzcd8faprQS9UbdUSp33ahdYLKaMnDmEErc2Q/MBcbFImoAq4TGJZzyJO5v+GnqA9T
sAN6f0r9wL2HUf8Nsn/S4UUog0ZTV39rZn0ukIkeyfkDxsSZacDYtPzBZafWuJBoAJnjoYgKkBZx
NaZi6Nu+S6jCamh5geNkFoWpaEq39l03PcrGlCHxqorGjQj/UiBfwVwFzg3lR2872KINSSW7X/kA
ec8idchvaeH5XCxvV1HD9IY+6aE0P7StjkNOtuR+lM7tBUwxX2qrwIj6oQxB8yVuv9xcxhQfBLrA
pS+2iTI4UHWbTuFWueRQ0jOZdD7P2s6kmzw/zA17U7ETzwn3rvLBiraGk0zS0AIAz6pio8mQryAE
kAXzW1rpCKwTmU3e64rL7pR5cWbdsk5kAzrJD458BUz0GKxQ4zb7ZiknigzAPRUq0uY9oEKhqvA7
GPE53DVcsu+MaCwgDprjKpIROv+zoDhexZbRugljwRPgk+EJaaHF6sCcRKU75dHqTbttfho/1LHN
PeQngh6/OtEQgyVbQerq2XD+MOXQKMvWfzjyJFIYcFB3pBazvhpOkEHyv6tszDVp8cgHQJGWDTFm
sVsb4cMyYNl6f3kS4BIo23xybrcu8NIr8WBZ6RqArQqetWZDrSjft0vtaMpaLRwVD0dB/7hjmYsI
GImPHxg0fQ2cfkbebhUCBcEvXj9cg6BsBWlAXiyhJiLw3SBl6pTNkgdbImsEdsnSef3p/fJWbc45
wFHa+i3GWKumO3eG56ZPwyDzyCXuH4WBbIOYd7YdZRveD81biqItEi3QeCfvfmyU4lqdlyk2pKBt
0Je4xN2OCPVzzNIk+X0BPSIDLEfCORQU6UG745fh5u1kERYS63JwqQMLC1Evx6w9g6O/xjC+TDEY
qgkNCE2l/I2JxPGn1DUkZmYw2P4PoEF6LpMLGRuqZKqrslYESTbEqt5t0phFWjfzwm3TogmMrJzI
Thp/GBKoffEtPZw1BZMw3fEVU9uX4NLaS9GqkK5guFOE733J3Cj/YuZ3SK8aMMo5W5yWt94pubyf
LELx+CtILC7nSHuvbfu4A2h0r5J4fzyQKZaXq0+6xc0tPHIy6YamS0/z1A8w1c4c4KzS0oPs6zNM
hdovWPJe+oUOV9Rf5ZIZCasdznkX5xkSiNOnuHFhh55NW3QZADheotl0STHKoousFGyVMmdIDU5H
nMCQML3n6RgIyZ4D1YzStp8wMxyWzxD738MbLO7qkfyJ1fw9PKh9l4UuYOeJAI7zoiH1CCbU3P8u
morSfuNcRAkv1+szCXqW+oIcEQSHyBmX7CuVAa5olcMicCKciBCxH9YDDFKK5dWbpfiHHG78uawX
bqf2k0ZQATLuJ3m9MX7tNEdEaiu+UOGxUvT1KHuDAFu1Ef0KHcGfBt6RKVc/lbBInUOgT355pJCw
OzHl7bzLinNlrkSPrdfXn1OiIFL/y7s+A3mYcWfGChB6+ZKr/rEVOBtC+m6Z70XugS3mPzvOBN/e
MbqO1XTUkG+sScZo2SBnwFg3fOgLAxTKVIDxHgKi2zaoehTs4njhjk1zJRX2cYCqF1fuPUyS5b12
JD31A42TCj/PrWO/07HhAAnBVfITuCZmhzSqcwm5XkcSBdVKqYUq9Yd8bcgaS9JhhhfliZK44wfJ
zmlSz1kEF5+44f7le1CO1Ts/3xvK84Xle9THJfK4KdtU8zMv7R90kQkhpZmjhryqFQdIGb7ps05j
Nk/eWBYgIjQB0bPajb0S6dxhjPn57y1gzyTQfIKywPFUq6WtVvvtyZvz2jxQkWW0cmAyLQGw1lw/
PPZ0ReoLlYZ/oonEiGAYOu4EroCj4u+qfAG+Y7tDCRGF/gQFomTBZ/Jazdol555yM73SEnVfFknt
LZTvp3OY1YbL4RKH7/tOFJbcGVTJNCwY8jdt3fIraXiAypAGjdMn/bdlckkbL14PqEnzTYLNnsfs
4flqjZoOrKFxuwsO7+3gqzaRN1zyZP2KIunQHcuM7Hs+Z7hviEOKSksbixvM27edXH2N1yCJcAr9
BTbC7LoRnWXirq/s5h8N0pHB7Ja5LBmoXnoSyeqPd7jtNUsuQbwooKr4PvmBtb7vpryW69LzA9Ey
y+bI/PxBhie/cc7i1Pp+NjJnf/jH/O6CoXcdoBeugXO5Ycq+mw5jNtXu+Iq20Q63uV1I3tevw73c
I8R6WRENrStmhDzE4McZGziRjvbwEHjtigY+WPPVlnN5mZbKQ/8kGV2TnuyMJZvp0qkNEklyBQoc
//EA57gj65WH+KPyNjGZ9MygxP16ezjA9sAVBEB4s9xOXjIobVzQ+L86ZEpoPNHeT298dKny2LbE
SbT1IkQSNy1XAHzbBO67Ommnofy2OsdIvMoSRpxwxFkrXIj3o5sLEt5+iEb9IS2jV/3Ljxdf9GAr
RvBCUNDvrMQcQQ2Rs1IOea7wZp5fNxWm6MvbgfNStGs8I2mTvc28ARIo9dLKk/NL/9CAbGvDL4Wm
XbV4qhEIMFHcsrfTTPIqoNgKIGht+unn+1M7evMDyOjnRMTrtp2sy5s2Y9wH5zeM/nkjsQXJzNwl
0ddypNKLlT6mIMSpK5z33znUfTHSGnqjN6c63OTFebKNBPjRmsbKgiuzn1S2GHjEjj8VnP5fuzc5
vo0Q4bB+Il6oA5r53arwU6hUJJgOl4QdE6F3cab6Jg9zpwTkl87jgC4bh9awQpNDF+ASxUUZ2dTU
pib0tC5H1RAaPeQtaaBL6WPh4/N/RgMTwrieOnVosY0jDeoDwPt7DhB1Q6H4vo/wtTwxOxxmW24Q
ooI8se6etlkcZiCcL5V+JZAOPPRJHVy9tcwL6T8IVQy66xGzfq+p3EVk7rVQkiQRhOUBXVPfSGqa
OANy3c+VVoq+4GE4XHfQgNFROtEO2htFZlmgLjuzTcd1sia2jDnGQCmQgE3yr0i29+VtUcpgw8E1
433jcJBFlaekKoFh0x2Q6oaZxzv6F75yWT5XWwD8V3n9wiwB35fyERxEIt+lCIUkIOfw77a3vAly
pcy5QjDZTKIvfH5f/RSfF4tuukuPsX++ivkLYggh+kKzNkqQ4XBVYS6C9cigV1QvVh5iOYjH2TYD
wKiduDs63I/MWt8wW7FSwQVHoZaUDZAMgeTpUezVlw+LRMRlQsibrcYByahnuykcSz5EKed8Iv/4
TKMSLKUPd8hga3kd9f4fQ64FEfU12LMyyo0YU+0mvITRX4KzaM1UwAeF8+YwZLvirPaDWX3XtS3Q
Yq6Cu1tvQ+R0dk7baq41jC/F00q+sSBCQemqVXThfBv1jO4DiRHTmsTCaKlumxXA7h+7mk6Hy8d0
4FjNocHVciWI03mVTmQjUagsn3OhNk+Xg/QNj+QQTeWql82w/wTf0PhOgoXkVYb/CrRUzKH+0om8
dP5MZNgwp1GL16sxnlkUFF3nVpWJfF59F7NAXA8aTMzhs+U6MiEBDl049e91cUsTOaLXCX0EjUHY
Su0PcSidv0IzjPuNw1RUiT5xra3Hd6seQb94x2pkirn6sXft8T/pr6ExnoXE99cyQs6u62AUCB1g
kSNeyw5G2wfSUaUmahIGOIzpbWFi2XppnxRyHEhfMM4uZM1ylBpo9prkLhaIshmiaw09jmlJTMKG
JCa1qIQz6p8HHY65wJVWDgPdGgk4yRZnWG4z06K/bwuJc8xmbuXuZ03oUI8JjrlBIXYbdEUkUajn
pCdPGk9hWkvWzq/XyvoAcVNAZSJcn2y19Ad2EyEqr0OM42hDJID1MR7XjQVLLGhKjLg7AI31EAAH
CRW47UjcJ0tpf+glqZD8u51a0xnOF2q0fXWYVpdTLn7pNEWIjp25EMrDsIBLnL4l7OP67eHsN1rn
65Tlbcl9l28UNOd4AZgm+2mf9UOQzaPxV1UayHxyfrWM8/Tmkx0W+owQOQUQUESWtaXWUvb0yXU0
vJtiCRLdQjyElSBfI1F7EsQwLeqZCglxEnmEz96Q7By/h1Shw3e5WV1T5VvhvEf2tlZRWcoa2u6t
8ZiGgkgav0pA1DiuBq6kh/fdYr7hakupWECzBFlkhcKU0fkxoT6pj3UFGaMxe2OkTQPj3Dg7laVF
plf3ZRfdQrFEC68bO9n1ylA7U3iPFmhUALkK6l1HXEcIeKzoDbnmb826drq1G9u86T8WpEbndCEc
mxr+hUxHbAMUhtBTLpvVoMr3DBKCKwJInu3o6mFnIEvQS1GQEXRO8hc+nUoeUOMuCfvhKCiyRSN6
g4p3vzQc/GH9wgCTuv9pku3h+HsDy70gPa42uQAR9NKbj6BniyUwzdDV+zSoGJO147RCxtwQYFqG
bt6mHuxNofhkriHw0gMniWTl1K0wLr46fg8FzO+NVsWYI1VyorIWQnP82aVrkhu7GUV3gryQa9Wh
lX/AEVXcmAhK8DfxR2daFjBn/oQsBJ7I6gmI2Cbmq9f1on8XaB1LlfYkHcS+n6xVUpcsixStH+ZR
K1+ppo9w4bkCyP0y22NI4ooQY0kAGm9wlGwFo+qMYhHom7ROkQuEyjYUhrdBOdkR5ASB1uCKtEqT
cftLO+Yw8TmGRbJAaDcqLHdTDA1EFRoyagGM544bKONNdPrw7b83V3tMTo9evVjPXyguinik9YIR
0nq8XxYvjcg8263ji6cl/dLSpSdBVmNhehQfztvfAAZpX8Kwh6iK2LeSQIi48NU+d/khy53d+mBb
lkWpHoro1IqRivh/E3iqDjp1DkgXtO3CX7RiK+I+YsNo4ghjgCGRBg7os+CwT9x/GOMuiR5FDqtJ
FCN4hwSiIvzsNTaf0qo4gkts+znVxrH8QNte/cf3Bm4K28EBpLLo1IIUCj4EFIlH+ISkIP5DRY7N
JWc23QnF51yqZg1evYhUuw1mi8Dzy6PeJAWgW+6hAWIQFn3ksPHBLjicycwtVItFZlZCzWzq4Fif
gVVccagMRTmJW7l/Uk53iuLImN1hFYQwN5gVbVGv6NkDVoTO5vEJcUurk3Zv5+B2RW9TW1QRZkYk
uu4fWm1xF5EZZ2Hn2QS1VMm8Kk45W3QbQDwklep6B7e1vs8HKufLeMU+gwSUyHqrUfGx6c16OWB8
pHf1Gzgmc1YbsS9qAMlmfpRebBliaIpz/C+8KymiPI5ezpb1+i08OXTYagBZb893PiAJmu+YdD70
kz8fFRQWuu2/nLMt8iD4eumEYFg1W6Myqsg8f91Ag5FpDTxIBG+LvRlcaaahMX1ouJBJt7j/fiO6
qm5sUqsmojAXRaeU6mmtfI11WDYsOB226TGNQcow1DHoQkp0PqdRTsGqLRciYBeuj7F99FkxZOGC
q/Ba8OpT4B+g2liV8jHYtHCxaAZBzzDzOlHGDXUR1DMU/ICi6OwEFFWWAqsg1bXiHO1j+8sPK8+Z
xO2CLt1SPjeOy9rZTK9PDfEH+NI/1dsfPtcwA/EBZwUjQz7odNwHGn5BZvyHzFPu1RPJMzz5BLHD
mS2jGQHmIkoxSdAPM4CAgXixm/vKzg6b+ayGxEbjqLJ81Hw1ovMs2lJDQMtXdFRjZqXVNPZiBSoa
tiqpysXRyCPvXQQ+f4sQrvLf32Es873WawjCYI7bKc3su5zXmBsA6oiU6Y/Gniku8Q+N+GUBXR+M
9/xJLLEfHe4Ygq227J7lbv6Byxo+4RsVPUvZiB9aFQLkRGGVKgrLdWNxSOmhPE3ZNnGL88NV4NNX
XxVG6A3YVf5m3I8uFQQAnw0/AF80lx0U+xGmv1ZdPzcd3NcH1kenmMpTX+2eWmdOS6iTsEE8sxt3
hhmjOySm3GkaR9VNLXDDw5Zq70RDZwGNYZhY0pbdREIY236gEZYT8Sg4W2ANm5p4zA2cZUTUoH4t
U5H8Q7nQPFzlKXxcNcdh/e6bwUzTkh+7ybJpxEDH4X7QP5TeH0o0YIspk7Vs2+dpxWZAnCAHeubl
tkd84w6MgQRu8dxJSVU206Pvi8BYS4eygBZQjusfIT5WUhlPGY8Y7WY/I1hvl1qQR2Xii82iW2Bs
4i4+/8WueE+WzBu2QzywNs+NwSCUwSVzQhaJbR88ZEWb5Rg/cMAtP8JUWM3DktuZN4hUtOTaBntl
rVkgl9vtg5Pn+0CwrhzRtaGK3Mhp/lXUOPDqL+wMtv04kCT2TRuB5+7Qz5x+pxGoNXpOmVVsFpXS
4+3H+1dBydKY05a6JELUfhNGVjImhh+3wLkkKZDzOV9ayo/eujTKHLZ9GAv9+DJu7mmS88MJUHVE
UWxedQDIYk02VWuPf52ZSgC6CZFR8A62xGXi4COXHUscwLWh7e31dEpRZwliOa4YKEEcH4WOJty/
FapswCIQDU0r/L1velwLWocOcpE6OybeTLEN+MOKchBCOJ8sw6gDQ0qCwCZl629M0Hx3m3DmoSPn
AOQYIOsJRnB86CTl89QMb8dg9pJ/Ww9EAiSd+WFQPt7ZqLb4eTwsXOeTNAhjWnh6uugHtbHVhZrD
jTRU0i05oM9XsoQ3n70OcM3iLXzYT964ozMTfxlen+yy3ZIevEkqr35XJ4/7Ekhg/vlQQP62Mxql
aihw3ocUXIHPkLcfr3XDizFfWw2gW5g2P20Yms6zVqSR9iIfHGWmyUOgY7ku454QwmPHGiorEb2B
7FQifxFTNXlV/pc3Rn8qnTHQR3VqgD5FJbsaXbLl3KNk8Mwb9QgXpc4x+UIeQH4zVOhjwim/Dic4
IIkehhsecdiKyV39WBq9OX+4XuYmBSbaQWQRTUfsqtBsyA9AagMCs8Icr3wRgnZVqEfDMYpCzw/E
GX5PeMgewnLnptPWCjX8xiS7p5elpVO3v2XdbQnmzen26x4kh29SsBuApedWsM/Y1wOtq6BiySLG
33axAasVwpywX378/TIEAaw9u7JCqSd1vx1YLLP8fbCCzEBHuZrfMsOD9UMDnI2ImMqSKKz2bv/U
woU00xwmrvJ5WCNiINmp+XEsUUVvVdXoP4yNNqiogwlR0AWBVTtIdU7N6hnUbRwYGRoV3+Oi3Pea
WROTGj5mdh07zvDqDIEdmM5YXR3VWEiQpavX6AMKxLL9z9N+ft+wLuUfeLxVJ8nAfDTFsKq3wckI
tsB2GEsR/M27Aikj2hcKTkXjLJkVs7M1L5OhUEaraA+Hr1b/MZJFNumxCRqx1cJRQ9Z2zsh3Q41x
LOc9Fj5WL/66QXlK94qN6yrPM3E2FkSWGSUlSVnG1FfjfOdkQLW1HSQdbKy7O0kygOPyn8tOwjia
6u3XBeUPrb1SM0ZxJHGNpATx8cks0Kr6NNdaj0EZMNScE4jEhRNemBDDI1H4KhMXWAACJO4jsZfL
xY6Oj2qVjpzw0praWiMAYMz5f4mYTcMiJwxwOQPPPPo9cyM/m1ljv8r1coLyUNE7Lxt7QPb/BxUB
3xsXK8X1nNvpwoZkfWm4L6pjmaslYYE29VCyWEvFr8haTHfS8/Dm3V0p5ex8XqgwqJqidZGOls3S
Y8SXtggVmEaait4C3frDZkEJ1yZuUsz1gm66QEa0+G6rIOvNAB7EjbbqUv7zSuWzP8bXGsUyJJb6
DaaJFERDI82v1HL0XQdXCfe5yvdiWvAlJCpg1OD/gILJYwT75ZOgt+LE11ztwww5NOl1Ep3M95ON
T6Rj0JXT5ROLLM/qkwkbJVp0RR9CflWqas8Gw61uXmNIMYPvTcXgb3f41MAbz1gq9EuzQSrWyMwO
JCq+/dFS+g7+g5vcrD5TSxvJsA3x5dFtNxYEieSMs55XwMp7l5WRToa4Q+d+AshIjphwn9QiJ/x3
WtkvSL/Sls/hYtjMEzShvZrdeBTjFbyp/C5Q53MGpoNEO0LNbl9KSzLhxQW32hw3jzP1plemTUat
0IcUPsnVOqhB/O3a/tVlylM6ZNLTVscWSP0lXiFEz0PhYUkdDZWonCKNvGV/HpYLZ/+9GW+G5Yn/
JbPSIWvJpy9VYVrJCHvVLPNZuYfMsiEHHR3jpNSnMJQ9XVRgFSIHkiLzpfXjkSTGYU7vv3oMceS+
puxT8D1DdtYTezQxauvgoi37U1HQwOu4TfoxpzfRyzou4mAKEcgjkiia/iucm2EZ/isYlRTyswKY
jOg1b6lkH9BSdsXcs1Cto6AlOBFfHSSXa4NvGU5jRBxhjMk0LRPZncgakh2fKHkjLKbAR3tuGWld
7RCDw37s5GxabROClL0wzoeG4gTMz4KuCPvzx2IB5pd8B8p3ogbGLtWaI0FimUcDIMguH6TPCc0Z
fwHakgcAgOTHoFCHVWNdc0EtceRXlqZAAbtOkv8R2EcXBtAX9xzrQKcvKJK0wnrYFkHUJtMP0UKa
/4bJVHmQPLvzCNx61flf97GOqpC6QP0UFnSvrY20lIrinDFHKAqc3cAeBWw9NNhQt4fc7KF543qo
zvlIlZWDLrgmioT70dTZxMbk6u/CJ404DKPUapEDqkIhIlXFLhGIaUMQADiJYt6SCTpEE2w+JraH
+4mb4ao7XbdJTQ/EAsL0J3WXpwt1NHpDDLdHvYINEAGvDTl9eBEXZajqxkSTugppRqV477A5Yz5C
m7Oj948zhDciIsRmd1B+eU7D/7ZCgiSTld7eOzeMj0VxNMhdIFCNWExa1QFtF+vaF9/wrNDsg/8l
v/OfFVDUC0HH9ZK+I2WRvLLfPBEAEc2AYlQquJogwgqhM0xiuSaJ5lh4xCX4W1Od1F+MXyT0iPy+
M9JJnEAgoiQO3rraxw0C+acw3qzne+X4pjechhgn4sle/IE5YYUFVyeO8Rf0BvLJJfUykN6KFbsw
J8cnP8076dfYFsRKDs6wDEjDGg+nBcRa9s+0i+Jr00bYYQsbJqTXZ3ciCcL7ffVZnak1p7Q5PV9h
VWFZTUoH+/Yk1BbKd88YCAjf92T9kqJ1C8RCRj7evKocsX4tCMeRa5nTm8GfElg4Uq9Xyx/0JZBG
SwDrJ4KhYQ3C5EQ7ATCqvJU2Msp8WN3XE6eAq/FpP5QNREJdrAOet9qjeaZSaOfv8lUJI91Ug5TR
OEpy5J2OuWfmwWSl8q9Ebiwed1ITbvdCP7c8fOGBHoTryMvXXZKphUV4+X+5WiTmaUSsFnQDpeLi
BnCYitlY6zKZN+5ka5B9sHN/SvtaLjLhBZ/8otOw1bn1a65PhvVHmxs5aAJk1vQdKV/C9xYt/M7s
fGec8QOvCXFOvT/LFjR7pE0TOKuvGZv1G4KYIZ2v5KzwS5/U55V7bpMY7SvNWRy1JkkNRi2vKANy
mLIW0kHLbsNUceFFEb1/vTtHgw97V3H7y02pJsA2blFew8T1b6sbu4axP9QkJVtWiaTGmFWSCrk/
v05JFi1Wtt0nrEy3NoEMpk1THGMK5OLGt9ZN7kI8tZesE0QK5HOani9Hm52//v0OFPmZf+C6NDp3
0krGb7JWvemnWwmjGjhv/gwnCdLKzZ0A0tmGtLd8mXeQNAT1blhbenL9SFI5VNWygl+dGb1oOTWh
m3IJHmtP1ktimhcZhfOtVhGC4f55DYXlZeRkm1Wtg9XQp/3wIlqMvROkBkRItCT/m4rea65s7/YX
Ao8udojzY/zu3pb2Z1CtNJAXXdlnHzwCmpq6fm+Ja/Y22KJzLv43g4+3UVg0MTulhO02gLdLT8pU
Ufrt2BILiNjU3D0frnAIXvenjfAWJOSwcoYP7A/3MDpYWFe5rQ59cvRREKNNlhvST2uBS2WiBxOm
gLr0v0OusFmcJXksHa7tyVXrH88BQBpaiRFvmGdlRkbYV+wy+fvL4JmTh4Jy3JheOvkha0COLyLO
Wu3BO1Efo28HSJ4atG5CjyWnzLE5cymv7TIv6yI3wmCP6bPElhlkuysoxT9Wc6YsC9r9fy4E0IeQ
GGxI4J6Zasy2la0Si0Kl4KCTUa5ZfN09azjkSXyJVmme6HJrSxgHh0W8/2s9kKOmOj4smHNkCWjQ
t4jHeoseNEfk6RGtHId2Frz68F0ZMLPAXc6ExJv57t33hyIpHUG518XBrl2249KdZikuvmBKUtWT
eC4OllF4/hyYaOqnbx4w8b2ttN4iBJwfXHRQdeZTcIBTSENPpnOtczzuzBzaC5RW/S3hbdiQTz2I
2bCQIV1sUUfA+QNaSRM0D+tpJDWVX7iCXpW3iUuc1Wuw8ikwwYLG7lGBdYnp7EjbV5SXQQP8b8L9
zt7kM8KJez4DTwL6Vausf2kyjb6K9cf1YmKlF1mZWIsDdb+RPzYmIvbAP+6UMCyekzP8AQkQUcSt
64nRgeR5K/hKaDiitz1gF27WxBBGHTsiO6kDkgClVYjUEvSQnZzJMxn+I7QtDoc5+5iWoJ6zt2sY
ZL1GdrguICptl/J23Ifvx5xFEr2IZZVrYaQbRNv55KD3zsZ9laRGuWDvNviwqDREEb2SkD76b9Vr
GwdT9WMYusO9QtcuiUwKTZ0b3iH4Mk+cJ2s5Va75RHnBjJG+tKmqLRb7eUmYpTAk6ykDSzuGyGbj
40ns+a7MC6afIkWWY1IDzaegKfSQnLbolxqTGtPF4X/5ZPQk3DBfl48pNLTHbGawHyIBT+4lVaNE
ZoaHNQz0A7eoHo5JdHFdjYoU1E8CrzIj3Yg5XRBjdR87ZcduklgIoOR6sqVPB0ZHO4ERCTp3HTx5
nqaJkrQAuAkBB6XD+BcG2rye4Gb91Tsczn23yLL2U9suJJNAdzWDiLkbA5couV9sNJ5gK5+J24g4
BQq2w2Litz+SO91tBM/qy4q4DEL0Erj0xCa52ylPemmhkIQPez3VsKp5oKHlLVLO5hVjDW1KFUM5
q3EmUeZizUa1r0kZErbG7AspPam8S0AN9ZiVbql70jXauR2QT8tfsfpGmuxhokDa8y3lYAR4hmXe
jGv5HmzyJ2iagzPPlp1jk6Lw2G+5tINrZPE+2KATd2s/EWAVJOxK6aTVKylyMJgQ99tJRK8uh0hl
L6GWtPO9+QWJ4sQwjKKcXVnOsLc65emct61LO/XLfhOvR6j20wI58rIGQhvPE34wbVij/9jS3iw4
q20reLmslygvffLsI1rww6jgBKixxq88RJtrLxLXM9C3YfjKAF9SnIo/w1ir/jWtiX2Wt/TcBCTq
ruC3hOjOf5VerswWIQPKETskO64IiApcurZ5/DaIgECNU142/JJVd+xbPNwNjnCr5WzPsaxvtCKh
HZRsZnvzSoBuTO1ZSMf98T4s0YzmiFIjlewC6P8cVXwDubH4rd/BNtQPOCRRgd8faEhKUVgM/1LI
9d77DLPaKTxPYAbhRtNVBJ3lSZYISOrisvzUbJNGESztNkCkGsRP5ZE05APKk4pIFLGR7fAvu4De
0o9RnOifoSK8SY+CIQxA5/ePt9hE0p5bZO5gqEeFzngNajauqmH7IE1hihdGg5JR/Jyk/5dOASlE
GAidc2HwIOIw7JgU2IEATKXUBWoYMcqIh6ucb+yNeFlGkcjYr/Dw8xpM2rzdjJHcW1c69E/l/5jz
4ocfhBKQB16rvMo132lfm7EZgmIqPOLbqyAjo82yzSwcZDbMO4MVggf4uXjgjWStLFHbNRwf2BtI
ZyjT8c+W2sxOIjnf7yE1pDIFmAZTx2P9XPAd6ob9jPWq9B0V0KorHzQitCtUiK8UzvGqGlBMit8d
GKM2T6//XzCydAsHglgNjSkEBRNxktikzWUZfcllh/JUYGn8+IQvQbe/hkXSFOKmxEh0bWH3MhQQ
OFnx2my/AZxwBxsqOvxmmkV4cJSVgh/aiOVTw1hA6KM7WwoWMqrMcifQmKN4QHBPoqD3ZYNCIzfM
pJsjZAs/vgfiVQNQSVfS/69lfDpmYAWMaPdKoVEGcDgzjd6C8X5cPPmlVlkO8KbDH9B6UIY9xxFm
K+mMKP6LWV7q7t/OlJJrJVSnGPDlY0SJiOJdK6gLnKoqXZEEjUaygeLj8K4pWZjZhCdt94mCFR3N
negGOlv0o90zbVHPyPkAv82IwPEHXtavclgn2NUpVy6sVcKIa4Cc/B8hqX91aZo3GdNDVbOY0jtd
M4YyH0cYmyV7bmcp1Ldv3dYAqNAtNHCYHKBlY/6J3CvlHYwj+yXqOmedohhsdRJpRcR4kChIKxA4
xWVRe6TMa9cHAbDmKwHWcii+cL57E7jsQtwGHrdOIkcd1C03EfJ1QsqTAPrrzP99rxzo9kcuexwL
BSgC2Tbweov1Cz3pxxUYOVXjkUN7r+XSP/tFWe4xLMFC8EoVQsEfMl+IhLC2m6wi3xKFkTsiXLwd
uArFh7IJQKY+6Pzj4Gw5AN/xNybN9f+GF3r8pPq/yRI+EPs2DAla4vvozXkF/xsqBkWzH/T6XZsB
eCKsKUG6tRq4DepuZAvSAGE+UU0cWEgW5y9+ZFZR63M=
`pragma protect end_protected
