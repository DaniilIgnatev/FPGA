// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tx79/rsHAvdJAnFogrpqqzmGZ4Yl6s/Ty8O2MANlTMx3dHD/LEZxJKQquktcff3ooZzzfz7fR26y
ZxQqa2W4LXXcsm0Y+e/vvUlR21dBtS64jAZxUeZW1zYy3QF/gG657JxXEJdH8TdmXzgJSy8952Mc
0enJJA9vTFicpSEYKXCfbIsDJcrtMaeS8Q30mSA7xdZzAJUyjP3dyMSwAT2p1PCYJz3BKRE0Vsnh
7uqdZM6EN3ZW2EMUaVasxL/n0q+DGpGS4kzKNudbO/2ib7jPdZzzLhM6vHB0MfgWVw1IAdoqkVl5
c7GlrKTR0y3p7tsuYZfg/wj2w4dfscIJe4yWDg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17280)
MraIweogSDVzy1eCcI/HzlkcBC4OELAek4YrS/hB1zHfyoKtE55deKK+VQ0Cj1amkHCqtkvt8zlb
vQktXt2VbN0mFtzp+Sym/Qg6j4cf9+eD4AwRhzbcSWDYYPam+vjkVoYys3rz0S0PYQbhiyNiu7nB
ZeOtFXp6p9CIa0z+70aXPDhGBXXuO2XehIJMbpsfUB8BTbfp522QQaeGshkXjiIEjiGURSQGS0rq
368ZFqkOwsq6z//UP4HEGBuzz4N4eI7fyBOckXn3xMXxFaYdHM/ymAniNAJNXsLYOZBCyK+LvfJK
6kwkLUxxbVSQNEMslBicRs7m13M0BUiTMDOzcBdNGIJRPVVSsmFWehmpCaJF21j2EgO/2H0EzW3Y
RElcTLJ8ZAihUc8zZFdMLA0YZYTzL2ujhMszuz1AcbBW34JU9QX+07z6cmXF9w4o1adxxYDJmQ0X
uoM3KgFypfNJNTm9xn17F9v55rclVia5r2MHBYmLwBPr6twjJcZr5yq8K3Nh9UBN/T7S6cK7l4hm
fj9FSl+QS1lL+x/h/vLBHTdsqMeRquYRbJKttXueU+xW54H2zh06gPq+Yf3uoVEKWiiQgLMZTq96
znjr+hIXyJwRYvGMQPfX7tyUhc7b9F3KG9+kswcHNbG1OI7Q/1iidf2lJ/0FI8pNYWm1gLL/xwM6
zgl/493wyhuxIBsAugUJaqhFLrYYhtvJz8W2hLCbOZg8NP54JxvoKwFFwUu+ZDOssEnf44aEFBkj
k9OV8nHRVKAlD+E1cOqNVOYKU2n5IgijTR0OW0yUsfyFSrO4IhM0l/XYQDuKnFjjfiIfijnGTrGF
oNvAgLKTd27Vyl4Z2rLegzjZbBlCcUWvABMqFTzb/Yj/CT5w0ryBRrhm/J1e+AKbHu0kq4uP/Mgb
MERr3DzQ0FfpoK+W7ymHTT/qu/qMRXyehLmevMqi0XYyW/uRwJos6XY1hTLpOaje9LrJ8C+tEXcc
1Sg5auyoTb4zhukTaIAkXb/117fKVqlZ6QBAiz+E6W62MT73Z08h9M2mQmtitK5u4dStuDscnq+E
qlzKWAEP6TBxwaWAqpEcnnodOyALxV+TgxC07frhzmUJ0l92jKkmfuw+TdlgNuItxhkz3ncSswqi
LhFm0dP+8tH6F0qRxP/AuCwg0yd0hHY+M72nGUKbhdedFjMy/ElWQrikklLTnGTS+zf/O4ayeZaO
MUyP3BxBqQZOw1fbtBhDTHdHp5w8qdDv0wH75YsOZLxv0douwFh7gdA070G4B7hjMCN3MkI13ghP
S+RmRYEYEEv+rymB9e2UxaEDwqpf+CzcZOsleI/TMXqyQ3ad1N0jS9sZgk6CV7bTgfJezhnIB87T
hhHUqWmTVL62aETWSJOC3mGzEGwQ+QEbvGDwWHLVgD+VIz3onVqYP2bLhr7y2PPWO1PHBlLYSykd
xI78/9tmVmuRwQBky6MyQS7dTEs/of+sMgTdjbwdvJCue0EsvASsm0g2Apyyf5pBtDWSvmmGoxoz
Z8ZsZ9zL+oNzvGI1FpDDreGXd284gMYS8a8RksnEu/EY6r/pzrLV74nOVT3dXdONkLRDmGlMx7T1
roXsBMIyZHMgivyPWvKREqiFu0eigI7N8ZtBxQVA9ZKaqvytcxAEPiVTH3n8AeOGxbqiLbCVuwNk
iXIWiPaK6ctPaHcAkuUAEplT7CKMOM0OQTYtwMh9fU9dCUau3Np8cqSJEaQPX4827Kj0LPyyx0wi
eoEPR7hwnpA4/k4J+4h5OZ7VOfNCR/o/VnJY3irrk84ZKafkJjxTX9CSA3SLFN68b+fU8w8hZPtY
tpoKrGOyCMOCAsY95WvYLpRPZ08Zb00ZBJ6t2IdvqVL3/Wnd6Y3BAvMHQZ6pQ0jbjUL6ET4xWw+s
P0BFWkcFtbkKNXqsEmns2PPTjY++06J7ENvcXW0NCIezkaOVx8msUeOEpVq10bJJpu4/4XL8JLaT
bVQozBopjy1MPgij+AKSduzOcbBmRR4jcb9Y7PgIZtqkf+I44dsS76q/L4HMbBXNuW0FGQTtQWpS
MN3KrqgOQs8QNh/1tNRoAN1VpWR+fgsimhXKAbDj/mOLsJxO3uPaL8A8aQTEAHR29xjUNAPx0XPX
SADK04KI6EEkOV3lWu8lFiNEZUzZeevK2tN9lKDK6tN70ArFuJIuf3DOa45ymd8v4X75OvSFkneY
CS9CleExgWMlc9x8NU9hoBTBwm5EgSQRsum/mtt2YTiuLutp8EbVFI3BYNI/jW039kw/McuELXlJ
nRVa/In7L2Qbs52yoUlJuIaHWq0Trg1x0iZSMyn9nH+sYlIQcHWHqIiBkYmbjqEqsSGZJaweWv+5
KA2cBzNAiRz5PKzgBaHuhvAQH39wI2HUVmu6ox8BwqpVplCqHX/rIqnHCLx8SXVdki1D+RobejRH
NwTFyDF68TyAPWSP6PGfObrixyJ3SxC7t2YmZooZp0iPtScl/QMwAGXQJi8DquDYcHwvKN6CQGqH
1yCie5Q97S0Bakknk9Xi8Ia2Hh4GFAQN9ygth0TZJhwfjbHpj/JG+WuSJ8O3pX0B2OCgR7VT4SDK
9EbbF/VDTWqoFb/Fq+nsS+/i/y0c7araB/Euu+8r4FNNuJ3FuHiLdlrSZmUgSFOzVuzkHcXAfoO+
9pwOGkM++KFaxnqkW+Dp5vD80pNIBAd1+bld8XLr0Ma7QpE1VdLWtw7259FkZLi38Zsyp37ISJG9
1iuQzPIrBTxniZ75M49DKdEndyGaoJUhsOac6axnPQa+RrtmsUAOsWVQa4nyCvKkanW7Byuhqvy6
lSgpSCX8vKRz5+LW8wwp8Q5xJYg9oxlfldT3VpXKijbuvmuBSkep5lA42UWVeTAt7Xkt47D5WcqD
xzbFBqLdgm6vhR9ZPYhZLVQmopzFzypzyQiYsdGaruTduEkcFXyBq0ZNeo9UQapjYwcdwwNbfOc4
hhS7wkIbqZAKpX6PNX3ZwIxXEnAw1Sug4zwGAN3F+hJTXKrATG5ZGjLTaMRRHahs96h7dnKNvUz9
wsGcWLLyhXZjcaddQsYSaTRz1v4roaNoGpVwiifYjJbqnFfFiR2zb/3XpYcNfldPmkrd74coi429
4A5Ek7KwmS+/xaCNhaCvDF7LzzYpbwoKnxljVycXWfHN+tj90XKbuCIrBlxw7wsiIIcYLmgoIl24
W1q8bynwp5gJRQEOWFn8WPSH62hrBzjw9N2kxibida6uR02DigVZ1JYfrVAkN9v5Pv6HFwArHe4D
HB240UlG56owE6KZjeqbK59a7bSK1lLHguF49nWmOWw/N+htlWddoG6lz+LGYcZTI1ljg2ju6w8D
2z/KwuIR6Hgl8yt1xH6L50W+LDwqJYC3ZI//k50Qb3u3IV6IEgkuMHF9pAMPytQBSZD73YrXokHy
+XkPmgyhBtNSUIpU+3Ny0N/Ob2oDOfKfDPqiOIC5vZWIfnne7IrR71jlUFMIlHlY3p/+xsDNbdz7
e1aab1WnUBWCxG5G0D5vqIpYJ766PBylcZ8zySQD4/L1Cpuay2EtaumJfRq9YUw5Uz/R7+yplVPn
pyXmEYSMlhCrK5ctDK6lDi7VwCRJUuAVLxBIQOxysVdeDayuO5nCdEFKXCi4K5dANO1zFIA6E7E2
Gvq2roE0KpyhiA4Qo+/aELY4jl70Gfq3cxPCBTFKHyrXnCv0INiWL2FRa9MPFTqSvzU3Ajk1dyIL
wkDl0JAWxG2zLAMoq2EtGuNMHpLLXd8xuP6wGw975b6yAgmz6e4gc2EAtVmEjmYBPJ8kF4Dfbr28
PO/BtPikgZz2TLQ9LIk5Oa2c4PElj1bKYBKdLOxuhm82AbqoQi4jvonpjFij3t+ABX0BVIciDhYX
lwUQBOWQjetX9DMTCCIbXCU7cIV9sx7TGbu80eNdNEuFODI7i40n0AxcPMQkVh7L2PXq9zBZXdif
3rmgTbkzgGqYURvgXGeTfo+wPxcQz7sxGwAZb53/Jxdkh89/8kyCzNlm3tYNtSIqIbZ3jbhX/5xv
Kpoh0It82C9zgSeKft9TWKA6/7RFRqHpvQvd+HNRv7JXDNV8KQ+bMS//zHMyCbrImwNPKPY0T/3C
enz1QnBUpRl1WJzGyzWmHVI1siAXRhpxmvLPsfsrs+gy8yPrkHuVUFnzJ47jNiSP1xENtDWu4kq3
oR55ddnw3NWzQMJFDaIibdyKLz8+ddF72AozWSssMpYCubFSqANA7eVE4OX9sJR0yI+Ff2Xv66if
x4fdthj+hp6fvGPNgSmc6/bbI+Nx3aakaJT9RDv1XqfIsviolC8IL8yb2hz1o1dj3Ej5yEG79fJT
elAtXoTsb0JnMkViK85JEWMTstuOSXVvFYE6NVkDJBI5EUzVfuvopkwHx+eMN9U3SFVnNsV891Fd
9Blq/JWpnbPmwkkJTqPBOSK+jfqc6XGzQqT3pSThR9NZFb+sM9Z3Epsl9zro3uvF16K3yJXNQMvV
6OGXvQxqMBBmTY23yIax3jy+sbUg2Vna6bYW+68mSj9/cg8EFXjEehIeDfq7Pf7qUMcT0MrMv+6n
kGvL3OU+X88hL2O/RFXS+aGlPvS7YI6eAeux4hi01GUaoNWW7SMAMHf8iH5l5Ea4EXE+PyfkgqK4
Z+JqE19PbyFcj+8PqrxOOFLlfnAUsciyIJeHj1L3AfGtBg0zSy1slG4nHZVfIfc+TA87U40vpXyW
WVn4MgoUQwcmoEXIFI5dP+CVU+aM1tlt6mCzfqF6WeQmPYKs2xGShJfTdz/ekJ/lme+3T7AP6VzA
l+CnHKLS231anLoSSzb2hMDoJ3yJ1ZL4ag+7h4uZHa8OCbRkTqHRjKSoytb/zXpIvuGo2FkFVpr8
yx8LKH/2gzZ1PZAfrKr1ZkasqWcjOvC97ZhPNsN/e1e1yqkzNUCIketC32PJEHYM3IDQYSwNYoFO
Uwbg/nwSUw3orSxpOLxNHJ5hkHydlFVKZjCZpCZqVpFRe4kZOeINUg//rLYDliIJB/wmdqhlDaaJ
sLFB2WASxjqvXxZBjWjA/V1vCCLmx7SbdEvT9e4Whipha88V/G4VbtBq0gtJ0Zrqnm/JMEeqUT4+
zf+Sq+c+d1llNBey13oHYvbf6pgLDaENtIgpQq0fllno+c5VAJWDHlgjta21SCiO2P+Lj3iCerKM
fn3iSIbV1auQevH0SbHYYzKIg7f82cvTdlolLRVaVP1qp9f0FppLdIQkEi/IT4mZayUM/cPjXpHM
r+CJddu2qaGu8EhDrnYbno5+hxCmenKrHV3a/z31rhOVLx7NcNpew9y0y+JQKp5ZawvnfZU9MBvB
csTWH6a0AuV1I4jUmHlYbo6HA3IYAhEvrtCYF49+/L575yEBbii2OBnJ+l8wnTS1Cf44MBn2Or4h
qZ81cqJCbUbDYoH03qiF/EIfEqqIWMQ0/l1MUVlAmk/lsBmlQpvA8bgtHVwp+bFIkZApY2YxSJl6
3V1bFChTPvI0Ay+242K+3YuZ9ihx481TORtg1zBqPZqEIJgj7v5ASwpOqiIb0mfvOnt+nQ6JkdPF
tjWZQAYwmOqGZr9y4Yt1ZmKrmq5ymXIvdv05j/FsMWIvI1zISCbHul0hzk1ZO8fJJW+iE2xHpEE5
Hed63bNL39c2Ql19/Oq50HNIxYnUrpPy7CuGZZYxOun8vU7+wQhfq/Kd/reE+qK8ilJnRdVr/ySG
1YdsOXZY2U0S0yowj4IlvaF5jdEfM5Lu2X3gdmmzKMaoq/nqp4APO8FYNKaj1w7JDgex6xxyu3xY
RyAL54Mt8r11JolQADpCdc03fTxavWKj29Ot85CvTi+uBDkmFKfC8nVliHjdMoDw/0INYUGBcNEQ
vxmGCBytXhwaH6/q0zJyDQWSz2fN8IPB0MPuhbG0VO9RZ4dLWoPOhorPIOqdpNAX9HajHMdMPZXZ
3rRlMEPKnTcmddKy+JGNxm0MIlWy7Hf/rO3KXV+Jrq2X+SLQgo7JaXgK0ef+fzgNnYxafcZV1jvq
PYJt4+LhkmFBAX6jfwAYlpGqko74XjuBpGJMVJwHBxtV5oATrRm34fTtSLLGNbpS2+9BuuknxU+/
SfXRGpniefRw/4YVYthlFGufAxGkVti+2tpQST4+BnYkHq62/aaylvjAjLx0wEJWiBAY0l4LFoV+
EVaOXFkSu+F3ueOsWFqd3p6FECg/uvucDFxrjMXly3PMeC6PGgCnvhW4JAgZZ8g4a+8l1MhUyLkQ
r7+JKTrM4dD/JhalJCKuMd+TL+cm2vXZSCaYU7KMDdT47/siDTGd3yzeulrCQzjSEiDkjJwWj+4Y
kENliW/jmmdBiGbP3NFB42pAtddfx0eRzB+9v/YYO2kOCTGRUy4FmHmaZJ/BMsm8XvRD4G9IgbX8
DNktklOCafeOTxqPM8SbCIeaYuYn6YEg4NYtkdlq5C5nVQKTFSNhRSEkGHeO+w6HfTuw5yIY7qs9
1wYtp/0WkZIv2RzQ8iYRnoeHIJ7uZ07YN+71ywGk/dGsmRWL6bOTNv8KG/xWIfRVaEGQvTWbB85T
vafd8JGHAbgNnQhNyRaEdyMAT21a7oeUFTtuOKJPxwIaj9PrLyRTNJVc11bu2fVF0LkuGaC9tu04
2pMEYWhDpNuT5AL4MQOpoO1G8wvzt9ui+x1DpZq98qE0boJUiFQ+Yx0UK4Atda7VZLzzxvC/ekfS
fHNYC80I6KTzixI/L6eN/JF389EQwpMiB5QWTFU5BuVMr3OV5aXBt2zTLsZCFUnGWV0p7lrX/9kM
9OnhXyjfGCZfwcqAXD5AzjqIxlVM/jpB19hUsKM4tLSeETGvXapFvtC39WaTh1iSTCaAKY6d91QE
cxvhsob8eFVsGjrQvlUtxH37HgegEdzsJbFgN/+FEp6z/Z9IITzX81rWUidvRKw1luY822Jbmn8/
uvigushKMt7b1bqAJgW1jlHoRGuC7zFLndcgXFhVklnYL5j5xK94cAbmYTrRRDP3P4q0GIqBsZor
2g+5NHFh8UzO3NlIOeOGNvbg9wZuaz8l8q9dkBxTjKqmNY+QUdbqM+StaoGHohEhpF4qlZPsY1uI
bMeeqUS7GimmVDhxw4y8mT9SsOil8F6IlmvOby7DCyvlHy3KQJmdLJvwuoERM4rfRcJdO+zemlJX
LR1Oaj+GivxNQVXnoLOufcdZ5tEQtR9qLGik6cM2aEYxreMh0460q/ZGiVGgbQUUBESQm5M4cMF4
owFYyvVNJhQlXOOvJRdBFOJUPyXgPM5HU3QHjR2V6D0/9S5Y0UeK5kQR9klqueOBD0t/OBpdjcKL
qPztTYodhFM1Ke1GQTSIJOevND3D262vooUnYO+SBbqe2L04HM7+sBCE0p+L5v/ZL9XvIyaHwAyY
eLCBVKQajg8+Ea8y3c/4Ie0EHIG5/kVCtOv3NboG+Rvu9uWGDojPZPVXEzGy9pziN7Unn7Tp6SWq
wtXY9/ZEaGNFjH3R+izraTQKcNALpvYcfQWtqfjI2+uGscIysOCAu4S3gfblrWLF+peLPyhm+Gor
mA7x0V0rlwb5Av3qNn2wQ9fb/yu+uxEXqFEKDZM8Hm9fGTan//E41BXI8gV0aRt1QA8dFPNSYU7r
YJz0/mANBVP3QUFfXhfAZBX39GWIjC09xKmskLqjiM5YEm8JQSZDTKvpGMGltUrejTppMq9KXvun
HSPawW5CGynjCT7tOJpJB/b/nkBHWmBJ9SbA1uiQC3X6GPOXJblMC7/jbXC1PmBUlUCeF3Aucz13
/FSZPks0qsNg1rAE59OaXfxdraJYTe/9PTwuJij1/v6nAJbv5aALdTbnBXOfF+kwM6y2JPZe/+jO
dNV/0oUM3YxTsDhpMqtf9EARcVXVFvO1irIpW5GcHYMArGJ7vKcHdOcKIHO6Miug8ALdkHGv6JlY
aDxjLCp+s8X8DpT2271l18qjgBZzNucP4MXY39MMJ5QH3Aq/LGYZgL8Z4Sxn/sBfvT/oexrXgyg5
AFgBcSKMcGZ9ulhdd6DjjkTWORAu7LSh4/XcNi222WhOuZE+8GSR0rRMZlZejyJ8wHczhHUexhmw
D6lHlyCBuzVoe2OGdYjgSQUY83zXA6k/MqVUogkA3HiFLAEbMvBKO3tANVK9SE5dTdNlZGLKTwXV
f0ZT6WDPYrws/TKqjMyftVRWsvDm/TR/MFKnsGNee3lwNm2uYcufZ+tXhAlno3qJpCSf94RNJZsm
OTu8ZkYl479y040lm5oEC7vYhSBfGPDx+ku2w3s04mTQXr0MQ00lZIWGJjDThFM7nWjq/YnGygor
J0mS4HJ2mVd/OYHtLgs7nsGKfH32cvJeDWcOjFu+zFoQcXK7N2dbx75mQT4lz0ZI1ng/dsirfkAh
AxCaEVyzN4FzU+7MJukKpkH8VeHTQCIfuNr15V1pqyQYXE0MeytFx5Y2t5qsTOIUTej1PsB04/7E
A4ucT+wPJaBDCCaehC3TQNKmKfJs502SMjPmZWGuYzRzRcSDHAZm2QnOYVYsVAP/z5Sd89cqlxG/
TytQD5ik/S17txD6QjeS+3DoNZcnh5EhYRIJNXVRVklozW6DVBQGbMhHX5o//hqt0KTk5JleOGiF
tVXYurqCk8Ccoj4rTVrvvBbXMlXDUelPbZVpvKCAL1mMm8ynQ2kNrOYaBLzCMlgdZ0xlzjgPUZX4
tf+/eDUAl1KahxhOOKA0jpnfPN8gMGqLvRGM6VgdHTbc6ZbUkrqOsrohjQwZ+85i+8l5ZBxgQQvc
DBDaFp7CsftecTzKzGNnRyQxiJGz8o+hda1jTRz0bHECLRmJPC3tHubtpI3BDEs1oj3GKAIRS1/E
CHj+csVMJgKffxa/lTWxEe5mDX1sIJrr273C1ElBXlN6vzP1eZb0PSgXwmfhcDhNieDAB1ArY8gd
NBmZ283wcxDSMI9kKfiSdtI6aNV0OMtpvnjHwr9PVkKIaQWxRpdvJYE5ZAxl3f+uatbjpeibBf+g
8nsgxTs3b+NF5QQ1xWxoqd0/Uf7xaxuHlQMqiHZVL1Rsm4u2cWaYe0vfVni0PaGlidKw6skI9Wug
B41guf3pfymJdfGDd356U197Kt2knTqhnMM0KEo99BGMUy3najlqVMZn/lEP9Uzmj6fw0bf3XlM6
OYON5YUjYKuWvy9RteBI1U6gBJxTt3rQUMiZ1kzvShMTWgG2STMqZmJu6Jv7ATd/rsCxrYvCusI2
/ULpG+rSqvtRUeDUj+WJxHt4ZJopSjk46IgCNFzLsgGsZTP4ZeZV2K3yHSUONvIuJBZJETjJlAHq
SlY6DSebLoKrEXwfANoO1jI1+uNdXvbQlo/L18P82uCuqk3ys+iqDOGz5B4cwQw0JgekiIUh4mBb
LvLfZB13xDPJfShkUs0gMuH0liWuqDYwaA3sDyTjO/pFwQHznzC/hVdvQ1n6D1F/cEEEyVV6opPE
1aNbXi65WWKPN/Nnrni1V1l6rPWfbHXrb9F/m0audECiS8YGeT9BDvfHNqEPJShSszKbPx2sER/+
Dp+7Cdv8bgZxa9H3eZqNE9ql/9KHGI7os7a+70EffTNjlyrgIHHGdEzRRo89QsnZ1s6PvurBE4z3
6qdoMG/X4AxxosEcEC0/+k7fEYZyI0nWWPTNjoQCLx4DNiuF0ExpXuTjv1AEXuIJb+ixIQ0NW8M8
DoxZ7lIYxWJeagnnDtZ90ofUBoFnwRmVCSlhFaJ3oMA/EnMJSCONzXN40wJgCEo+dvqy7cISjKyc
fLWC58qAvsHze+APJsCKDiczj1/DM+rSolJxZC4eV74t7HEeQ5+qeQ9Zh5K9aSOywTaaELc9ScCZ
wLx7uH59A3m2ayV5kLVP6csnWNNjWNUtgZ4JPzDAy6vJbih/STAdYCbXxT1y53faNdtkMboLuAoe
N//jROWbtsYiLn9sWxOukO+Ltb98jUThwsoQrS/Shxri6RVNtgOLYWHgMBvXhHBcGMbSUAPZRmF9
wpmgQA49+CurBnKv5BFJK4Lkb0NmKINiNpCVPxr0rgJD4PDygrdrcWemR18uKmPZRC8h+yCE9RB8
x8oRXJ5xt/R08ah33Rmv8VE7KlKq56SUa2GHZZ9qYyoHFvY+tWnsVYWSRYQccH7ZrzJnKN+4Xkj3
vdF81T3Uxyk/5ljRD2HOxhE+adKjn63K+6C/4APOX607LH7Z3u2R03nGJjfZH2WSgB9GoPaXPKVj
87ftCbcT7KvxqIVv9XeobOV0rUWOXjGxOVbANoMLSR+0hd4kd/dFOLF/VIWuFsGauwdNYhaqMAXR
oNEHuN3wpAtcSigqgB74m4klNSGwZLA7MB98wNNqUSfZhJCry/kShDo/I6JfLshpMY+fjCKw64FO
qYkksTQrHhUjPNHSAni1iJ5Woc1c39Mso/RMlhWcn2RTS09EXufDqN0/D0bLDgvmnQnBg7D/O/QZ
KzVnSNeKKGyBdl5ok1rI1Mom6kiFhiONmzuypSaq468tPYEVOpsclDpDl6yhxP2HK/C7oJ21zWR2
OH5ghYgAF0kS4J3O5a6a+Emjhj6v6+W98tlwpBH52prhltUImtyEG4et/0H3dMZ0Gz1sVlx/5xo8
7rxnQC7JqnAAraRFMHOhCSnX+lnxVX0ATYn0xSB9+NFkwbawng6DhsuBO1uQyafvB3Lyt5kQoF7t
1IRWHbf/Kyod1WHUkp0E/E1+mTlXdPKwQlO3kRWOBfeqS7M9n9XtkbdGJICfEijXYccDN/8YqQVH
NTltEL5n1esclYD8QplI5aaG+9Z0AfCaY2qDw40lUNCeooC1DrZclBgi0a0H+2fh8wIr09VC8+ix
R7g94huUoOd3KJoVoggQvPhJLknx9hDkP3Qs0zBLRa2Z72MzEQS0uYtglxkujIMDV0LZlUNimHwh
dl7CSEUqSIl44gwY0RpwQETsirTjOlTi1XgpbZTswXh1ZHiF4g7pwkkWMJLS20fvDORQ936smfSU
+dhue8JIkE/VWzc89Rv+dPfPdOCbUZO4l7Uf/6/sdA7pb36bGP3HO53uHX3RDXTvwO5D20b/Z1KY
r2bQA/+Zpj2Ly04W88qnBKdLffQ/f1bHoflLN1MbnbXxa2zpAmonU1v3GsIK5R+ppt8Kl0UdyMFB
7DB3eVkpkUEjTg1jvdo/Xx3m6ibLwa2U4fF08nzwftyuNYUFWfEXsrtP868T/s9fgL90JCcykW+t
fFo6PSIWMnvZHqJGZsTKBjpE9mClNLTYDc0xgTEz0TY70jvuvhlrESTRpNWMC/HqNj1oQVAiYfna
DqyHmwhJMMGcVq9HY/594YHF5BkM/sdtVfT5SvM+QktSeA4gDgv9BW3576wA0veVJc8fMfpszLUl
oeQk1g2ow7IS16CFEDGn4Q3lwH0lCZNnj2ede7osZcoLkHp75J33Mab2UMSxYwJK+YE5TLqgFtnG
ub40Tb2M95eGwGzdsPw+kexd6yHF8V3up4sug1NZ+ONhAW9u/3IvT3OnA3FLSZQV0jqXbZEpVq5F
3N16zBQJh1BXLtVxvu5Ybt+jLNTe/ekI3KaXKir3mizwnPJLbvNamXQtMNBkVfAbluvnNZVxOoRh
QB2/zLZ8U6nPVmgl60/q1jF71CPYYVSXnEWBYJT0zNg2BnuIlB9UcBIjxzMMusof6WSluiaUxmmM
UqasKvOAfLO/gdpDL9rNlaGspsjHuP5cI0o9Gx58jbfISQ2kvE830JaXkuXh7m466ntNeTLNxwNI
Qt3Ren5w3dO9sQ5hHtrnkaIsJwRBrQToEtXX6+EONYHY3CzW2OIfdwRsY5i3daqQE7CPoY80PpUY
PZR/51h3VSmvDUqW32R0BfMxBkcNSmOotxD/K1InHWoMnz84JjvnCnZN/qXhDVh7EcVpXSo10Kp6
OF+f5UdwbGU9K80sNiIB1rbIeCtQhhaEd/T5ULi15+EHZGNAh+cVZoxX8J0HuG9yDoy1Qri0UmqK
5Rac0sl08hGJugM/5n9+v6B1S6eT3vLG1/F+rIQIHnTcMUvJKKwdWFbHoAutBW9BGGHhCUAzjwEZ
4uC6sUyGT+PA1XCHVc9Q1D2MMUFF7+3mFZwBLbQ+pEWC12iKCwDFi1dkx8b9BysmasZOgIrqSHdT
9rAA89T33h18LsG2jSjZmCcMynYB7JY8rX6sRIhPoiU1qyRSWid9rS4AG6sk2r/MfOhNLsiAwFf2
8vVWg3OoY+0WLNFs4kkZ6BpG9Yak8bL94SATFIsMPLeXPBYN4dyzbAhq0u2yohbpiACGg175P19X
3+BmGZvt4Am9O/wjuyK0fb9Uf6AxwZdyrO0iUG+MHHHneKCstntaBNLE8DuXqRZkEZDDgUXztLvK
KrtWDcuZgFK8SS3CJ9j5+gjiNQ1B/Gc4NgEMiiZcQmzUjz0OzAP8C7mAYEjd77unkSzt6/3SR8C2
z2Sm6Xv4atABuRZpHswxJQWQigX7pOxUaipwPe34KiqYegQTy5vca3PFSocQMvsG6xctF+24ebou
K+uj0IhvZkpqFCrypIWZifrw/CsZV1Q9Pr7Gqy8jsPLewpGUKUNyZ3KjdGmAwLQZWjMhrCIUVc6H
7sGfXUt0847L9WjaboTCwhYwK64cHTQhSLz6HUKjyvq42E6PMZJVlW9pDPkANzcKZaMrfYk77s5n
6cicODRv56t4yl2vTCn580aS61/4m5X6g7pXDGf39RUcVkhnV4BzqQwO76V02B2USFcyuJjK5mCC
KNOKXU//o5JBCsndBuCk0Pat4WaEccJp4N5RX4GjRp8TI3bnaBDU0oO6r6rR+oAi/mZBY+Y4z/NP
xA7VSsltx2JnmlsylqcDTdbP7pEXMpfEK2A7ZHuWLou/U+GYSGEJIfWaVZDzK1wm8s06K8Yqgz89
6ubvVHhhFtmIU8SibFxnihk+HihXMwTLvJCO8zXPPHYEovrP2VvnGH5O4ifIXCigC3DiP6PdVJ5z
OUYq83RVoc0yhJbisvkZG+lIKRwBXPdAvgwSZtlBcs4U+SP9BnRuMnKhDYLi2QtspFOYV624DSJ9
qECDmf63p5jSVxWLRXBeIWD9JuydQ2bDqzdhEmX1Om8+lR7JJ51wAeGyfXA33MowRq/i5eTApwjn
Lz746V/ODHrvGNevCfaOeYglUl/bA9Xu/IR+Gyza8G1wUOx7U2ki+rhRzKalSD6J+3Yjkt/eU7MI
olV+72SvSqoH4cUfB8w4wKrgMY8A01xRJbeNQ2QS2nKuIBDqR/mxziemp7aNyq761vC+24kCT8i+
vZ7Hih7fp8oo0QIx6ddvUp9O/GMTLDzL7S1PMFxLN52BGnpjCuFEuq3VgrCZxZJLHSl6oyfVMeBU
PtBly0y83B7g5h2/SrNPw6xRlrLxbxEwpFA10hCAcJlcee/n/kzF7cBJckGcDg/ovIuXqiQi5XPF
Ibkllj2WnPF0TmlrtntUsjCziTsrJzwACNyyRoUkZFuDb24Gu2Jarl4fTOF2/VXbt6EcDoQxZnqD
RTXGkQ9dx0QHqXUopP0SktZxOjK115gzKx/+DZA8GUvDaBPC4HKgl0ypVPU9aNe4IJTmFg7udQkk
21aYyFQQgLY0WXgBJ63NMgZW2h8bKIwxuyhCycKbGBcJOVLU0LpCflarUSuEMCu5ctkYHvtfUy5/
MIHUJLOCHuphLl9ueum55Pfr+IYGSVcYzMjpRN8kLTs4E7iVNhQC7SZW5NOBLPPw+VtoZP5cJqwk
SaMvAUYEIP3FQG18kwcK5DxApbeURa/y+KFZTIocPen010+w4OxO3Sl6Kp9sEWzk7oaq91CwJ5ZV
3HPhfNA1zrN0Uxn+5PU3qxDYKC+B+47qfz2jcfkR33FxRz8KDWCHcDVfRLVvHhxVqc6h2W2xGHdj
ygDz+2ykFQ3czc5CfQIUIkvS5jcIn7I0QMC48CKYJFTw9lqeaA5Rxr0jrjSAJ3+aMFwzyJUb5PF/
rbBlEc4vdqYFykORSE9LdQfRc7Z5IaHHW1z2xmATWKsjToaTpLxaieyXvuY0WdlcoBGtpcGH0ZhU
iJS4zNvKoCyZbateG59TF6gzqi35De+0RX5/7feHK7OZZZoyH7O/o0dbjVO4n7ZC4Unl3cYvbksa
gkc/pUOC69wyff9AoE9fYdNWRMzXS3IXJkuVpimHJtW46QEWWIVVTEVJNwcMWV4KoWM54NCgdyYR
Rv7DObJxuj7mTo5RA9Z8IPFMjQzzV6HYzyJLMIs3JM7viX4RI00gKILJ2f9sobmCp2+975oSDjEz
Rlz3AA2g6DRqvqjUlGB+SeXz9AEHZOyxFcA6zYI2Brhoc4CpvPT9v0TzmV1CSi6xZszEZ/XZ0FHm
l2z/igtw3O6bShPi5N1O92BMFMEL8oEgRNIya8Z9NZJ/a6RJmIb35hfjs3TKX5SzP+lhM1k61xkU
h4zCQu+pcQKx/+raqrZUHnQP7L/TLoWznxcb/IVBff6c9nTGsDE3jl4meMsCQMZuY/aWbIpkXBkR
d7kmcPnLyTwWrrtpjh6UmanJ6RJVMrXYETc2YuX6iIDHdqCd4bKqiJcBmNZO7ayUFrXmuaLB9vzI
cIomc0tJNTo9oQktgwV5RuP/9JkFd9ap9ysKVv5aBt0jIs8P5LIlHTK7BM/fqP+zImb/Cg8UaQtp
Lo9iZgK1g/obVx98vMEBc9HA9Pp5qFytFg0kqvfXCSJ80uF6bml1kuIcGtQo0/z4DE8QzC0WOUjm
upLvZ2ZRU7SiwvpZbAsmRKxLEKxhyeN/uMQAebneiJ/wFT9F/2oAl1uMiCHNsJffMVKWHrgUE1GS
p/ypMk0Icmk6SY8aFnIzI2Gg8/VsTTVEctbC+9IiFVQFj/vCaDiXNhKEi+8LpOIjuXytMJrtPG3L
6TCChTGLWaPckTEEZ9vGbFAy2OUa35vtalKwzjjFtYJTlIHp19Utw83T1w0CF+Mt6GYJ/tePcaej
UuerA4WVXK/Xav06OjjnPP4mbsVPssMOW8FbS9Wo4DCKD1RDps2v4lGxWJLybDSF/3YV47tabKNa
HsHYdcfkhob+kkoOKtdkxyWemtupCgQPvdw2vXzLFFSZ43LEjmHxbw6xQeVTvcCC6HF7LdOVAEnY
oUjhArBcJo0D98nSinf5ewJCQZfaS2ugtwLu2U0HiYpKZfd6Fc+4IdtRqfX5lJTPWbSDFiO8QNw/
ndjo7lhXPpntN/b4IB6d7pevuW+RooUIgKnQmhawRJpYvzLT9SRooodz5cy24FzQjoOWwR/Lg5bD
gqzruY23C1XteaJnR7gEEpM3mTQd6vCzHmAMlvNKlxxpOlo+DsAR/EZInFISOoaJPevKSrl+Qtfq
hU1q3zoio0e96nnhveIJu9ezDiFuPHFaXKDXcA3IG2Npdcc6/hkwJr4YjJ14i33+dMvEMLc1N1Ty
BVKkbzMfV+y4p6xBjqxK8mct74ETH9b0ApsRvCxhtzc1N7zAQZ0dVc6jpBv+9SHGvNpwrLT23/Lv
DuUeX7P9tJm47Oyw+Fslq34sCEOBPFHCtgmu5vmr9xktelyd7Lg+ZT2caWaS5o54kPeL7reOYB0E
4AMXhj/iJ/Ljcr7dmAwvf5ISXseW/4WLOWoKkyr0SOT64zn1/LxzNPbPNfPBmU3mwmnbpxQjq78Y
QgtRODilZr7ylsoASNijqek+VxjHBU8TEBvaKpRKf+8uROO9Rhc6yj2jij6Z0ptRQFh5MYvPuXsY
kE452Z0bCYvuGy/Nxessq2ij4emuknv3PgwNDAyK0p8LQ7Z+0+cm3rq4NtB8eXteMGzp3GVRnvBq
oYuNYHihBOKT9wXcHvCAqoUP8wevela+mEjjj8Q8GfhgWC/6DyuDeKigJQSm5aSY6pZGVGOYi7L6
GRce6O/UjXPtfhBVRfuaL2rh5laBifW/Ewh6SOaIAu4YMWogMQPgEpc8nE99M6BaWAMaZUiUJnxh
QUaU2prV/XGT2AsKVA1uQfZIeM049PHmPiVyPix9jdTsvm6FdDax02cVw12te57UCnX2PQQcueQh
O73dTv37Hd7ubRiFl1VCF+/fHXX8eYINTOHQLU8ICzBXaWvJjIF7UtTE+lpxJjSsjCyAVjg2ZSG/
mYDWq21ycginj9r5zvzBbdyitXTrGbffUwV45PUdJKbvyUwxGEX+x/q6L50xyJ5xieOJRQGkGQ4A
bBAyCrsVXoKj8oDiYyCZQrdIgSqt0d8KE4+Cq/0pI/Bili1KQrBDIFItHzce49SjlhWjcOoHNi/P
9OU2AcwRpIyLppgpdPeFw3DH86hDHvrz1kriNO1TK2r8YW4lGOWIVou8ve6FnTxHXs9+dpZMChLQ
vlxl1euhXFTQyMNisXf1GYKTbdGj/MgqTEvGtYuq4lYzSNfb7gquT5RBm7+Uq+4KX76CjQIauMZ3
E/Ds3XyBB1JB+p4KuF9FINzLLC/7RhdGS2jpTvESXXej+jVCDlM0fldG1xPBO+bEhNnBIhl1orUu
r3J7a8pMMxb66J/8/Ak3gHQyybaQmR6H741sKYI5ITA/Hgxjqr7DypQwFa8AGDjVrHWzK30PZ5df
9oaVDHraENHh2CBroESR7PTtIqTof1de4cqnBJHAd3GcZQRxDxSXzvSkwRo+tCmokr1MkbYa01HM
EM4+ASxqzAL7joPpQLh+1P/mxWldByTTsLcoMZXiAN7RMO0PnrBws0hc2AYCuNC2TScGoc3qMmI7
Et02vV/FY3q9KLLihckmDxmX1jDPVf9w2mXwOrvufWb5BKOOf/1tL0YXArziTfM8uomI6c5Zly9N
PiPrXCdn+wUmOLUSgj8IE+99PxaNmgzwWKQaVMUUqhwj6aTeGlBuWN1CMzpLjL++Pt1gG2ZyyKEF
2lJpjIV+TPJDTx0FI0zEb7E5kS+JaGFxbABIjfLjwbVOksymGq1lSefFB2lP0BkXvazr+yJd+vQi
1lov8JeDUxuHNdScCJFIdJAK98n2gQA02FzAtXuwqduYgeaCdfRijtw88NPUVeRGKw8jwWCC/2Sm
upGafYl4e2DjtWc1ChROhQ6WGWheYB9USwFdO+gBx1riCf7oWSoC+/qXKVdkNqk3G6jONhWbuysH
n2YSFPY/V1Hyh5cmeqpvUlqQ9HkfgyS8GVPh6FgCghJWHvRbi91Ls4TOY7f2/kACKrt14c1na1uh
lrAoWr8wLR9IKF52QzhOG2jDhkwSpEbj5V2I5nGO/uCrin/zVftsaIYiy3LCm9Yc0PgFtbMkqYnF
Q9xhbhBFykFm2aV/ZmhWChE3ynp9fb3RKK/ZdcQCi+KWxhC2fJy9VoQwxvilgGdTOBaZXi/IUW9t
5WurZmoHDtqLMHrIx5z7VHvi4wC2k8SxptfUcDkzXHvKf7WSPhdjv623j/E0WQt/nnnAbfwmiFrr
YeEvdq6/g4D+bEwaLsH78QA6hMWFxR+EsRen0cX8HsPvwPy+CHCG+1re+moROsXoi34NPknXY/4y
1lMBgtXhiztV/FXM8za9qtKRF0qdum60WDA2s5d4bLzrv7UGyUwmwRYU3adByGfs3jedUEYvJ3eQ
9Jun7hMk52b6NWD2eobuMndl3DgMX4ar7XUWad3qaxyqhT2y85wMARR4bJOOarX8nsGOlNqRL3N7
MPqYWdQP2lXV6lpGRkSVdxTd2bAFtlUbnxwYC58YAQ7YmIGa3vOuYbfDQpIc5aTaGclnR9B6mZQd
pjWZ/gIWE5/dl7av/UJXz0QtgcJSwAoFnc5vtXWvmuWA9kyX7FEZ4gd/AnhynK2ApQDI+uNj4r+6
6EI/TXpr/rliTvfdcrb55/dDHirb1I4oz8woIOajXLyc+mgWRQ2PhTpEw+i4J7HHn/mGEGLJrfeF
b5ChCIqRqcISUyxWYUkTWDCdC9ObN/hlI6cvuYYVCqez70zsLwAcG9ieKyjIqAk7NGYPdg5gedsR
+8fmTLcfWK4bPXPV4XegqQLWqLDjbjKPUG546hh9reHH7Tc+X+kMgBWDRkHp9KU9BYZgJZWn6ZWd
9aNugCe3Cw3JE+AFCSPOGJFo3mJ9Uw1dQkH3bLUy052pkRqb+o4pxZwnpoQyaDKOFh5um7PYnLmV
Z60VgiYuaTj39nOFu+sZ0R+Fp6FtVdVvnjRXfZRn3e28WUKqQrca8pMBpy4HUHZ6HMF814Q57hzs
yUjyg10q5IOh8KXfDLfzhp3MZ+DPCp+fnBPjh44ycqrYo2ZtLwGffntX4jByytF6e9fpDZiLD2ub
G87eR0BdTLNmtD5+PlaypmLxZA7ahv/4Tz0duH+p0R2gRe2Th0DqjTiA654A/kElBT1fxsoE++wI
hr7mz4aqq28uVtEkp8w4AuPdTSuRM0vTeNdsD8Pr1jywAHpJGJe4OGomoBZd7lMTTjj2RaseYsoD
mGfhoWk/y6Lo5kM4+gmkJfCTHv+cRfbNy9nHt6EY7cO+Y3cPAPscAUJVaRSkghKYRBL4h/O/VrXB
8TjnB8YIXZNCJJdlTrYiwTOD3vrDg5DgQuolILBHGRLiCTPHajdK9SHaCePZxZKj8pClPLVjFPS1
UCreDoLbCCR/1kUUQYPFcVGp8ff9wgK0T5ZTzAnrG4Rf9y62Az0RBXOfo/ShBAhUhltGK/XyHKu6
5godMNR0Zo4TTXNdYMYtEWTVANQp6sXCUnv5mhxzHJvK55tZAdSCBBhunBeBebGToJdeJ27X1sEX
PQjtZeF+85l/G2FiMRPQ7bxqd17cmr92XgSLd2P8VjBb3oKt+xqUl1Mjulq+fXS9NfJ4xPvGu4yx
5yaVxQkSRDzfbD7d++x+Qv9JM0kFLB1VSDbrbw6062Y/FtEmrzKuU6BxWbjsANGgnqvm7xOeeU+m
AeDcJqD6ut6KV61Is7aQGaTwiC9kEuYgco6/9mOAp4Sagd2v7JE2nOEBwe8EFN0bFakYS1u/Xhsl
8P+eciUTE6U6cwAXYfg18tHFl5qECoMQlNuJqLPvPjduqVNjvx5vNJXUR1dt0SuvLOm/lG1vKbkp
xZ0dw9+HUumil3sNUdaZEfC8Q+roiMKkORX8qZQf6Il3ryxzlWHsR/5VGLp6/BK0OyPGOiCGGSvZ
rLEp1wBJYdnSosFbJmwA3pIix3YQ4ilkAC1Z1u6LMglYbtGBNjkoqrZu+PK+6VezPeTt6KScumf9
4zNexGnpvCCP0Cl85sCyIbXhUCllKColeVfzMjMsed9skNG5SZudqvQXVMr0sQx4WtLU1J9Z8LTk
+UzxYzy8Fx16JvLaXOfxatzULZXdjkDw+3K9GaNGhngO0EuxgZIO5Y5o7YAFg5XrhBWrrPKjLc1t
bB3lC2XR9oGK7XL2ymIZHow5H8qShav+PSMP5XSO0mILmKgC41XFFTC/BArBzlhO1r7TZTCzbczp
WXTS0Mm4lPdjwDvY7KYwzWuyEXLPVicL2C8LbOhmFrSQtlNTwvCo4iQd3TTNipZXpKB1tPF/6VBa
O/Kdow2SxtolxsvRicLgnaacg81jb/pX4Cfcw5i72gTdyWz8AtjciI2jaWdHe0D7XUI5XurBQL+b
cC5T6W0rGr8GnDDRa4RKbhd/BFV/IyuGauRrH9hTIJLsrymYM8BdQ2nfP6b7uHyt9jD19t777tXJ
Am6vDh3eCvi/WILaLTL19eFaT8oP5HcOJ1el5Jlf2RtgBYkWtT3rO+cyVrU4h0PvqaWILTQKdjjF
ppBfOyeFY7bKBnxXA7A1+SdZJl2MfXXb1Xo0qOfLq3dp6blccuMmLK2icIyCGvr7x471dEm88d9N
K90s343Ulkwe0jHLi20k1OdZmEaoxdeAVXlZ2U1dkBES8+PN4zGEobRgw0ojbcDg2nv3X19uzhgc
fBmKXEBfnBX/ETnSElUL4NVW3sSciV9qH0f1bkvLHcfbVrMY3djNmmjHClDiZEtuREWTAxSJSJns
vfSyNGO+8TLEWXeerVf1E8rKNalERWtDuAXfFBNCvWZcaNcCTbB60/4rBhCKCcuT3kBBzIDXWeQc
j1w+2k3aysBxtkHvsO9brBkQH6ov1C12i4IOiqjKX/Jdr/889clMDwvKHuI+vGCYWlUVBi3zOHEQ
UBdtyHion/Ikh1+/fe4OP2vp9zuMxkGMQHHeZ30Pvhj359bJQ6AXnr/H4dFmzx+D1bbCeGKOqJIM
Y35hewSPyWRyggEeOg7stfkGGUgywoBpsLtFaccFAd7ZVnqV4kq1Tdaz/oRZIUEVBQabob3/zWtK
Mbju3+LJV9rGFhqns19L8d+ih8GNKwYyRwqLA2k8O9R+f4/3WF/mJC8YA1S8vsaWSTjLrtBI8oO3
69AgHQHXba6bOapKZYwM3u0TK650BRLf3i5y1avVFA11k+Thl7ShpSYIm7u7omeVRoL1VhNM+qIm
NGMRFeDLAMhTBbfXnjnkBKYusKw3x3lZxZprnLLrlv4X6RKxiRhaHTzsQwis7ylySraJyAwdh/DN
anEl0CHYV7VSCdIeSqeJ/2vA014cNLOxuwykuknolvZeyKY0VXSpAHx8TJKwpFHB0D4VflAcFfc6
AVUwZGp92o059GOGwttd6Qpjr/XoXlTGYTjAlHCOZ7rAy+hJlAagWcTzqb57NAeVtN8M/7+DIb4H
FuT/c+Pv8bIvh/PG4AFCBWJwmqj8VpmcYwHTEgDDOzz982OAxW2Ft6CSDOKPBcMDuE07R4N6e3K4
0lzoSzH6sLlRS91TUpTdobHQ0QABxgLFqvhFR2GcGsFGJKOSD7Md1Ge9HsJdy3/uEqJa7AJKb+lU
0CNjD/GbV9352xS3SP2HQFZXIRGRARivbBV6D1zARrbtRPKWw5VWRMtJEAEYThN9DQSd64l4rNMc
/XQZFOGRPzcv4gDvHxw8TyvGlZiBRTLZy4wLJ6h5c5ir4xvZiPTwGDrY4Ki0Em7SmLpOvSQpf9fh
2cBL33uW/64Z1fhuk2dlUMiyyuaWCHF7DuJA1Zc6eI8t5q5c56zSlNhqRXQ4RQ6wfbM05cRGm0JF
fLPBbTCGSkQpzitLUcV2RJbK0atuevtsToVnqHa5VZRkgoLIGIAEEuLwxJnDTazINsZ5YNetqio3
Ma+zlSzoGzy2xkoiUr4/GfXXP1h6jBggrsQTMc/+x2pzV/2JZqlQ+o6ip7VS9sL1QnOXL45uhGwT
vkdf94WJBl9HMJ45B1u/P+XOV3CZg/+px16S/rtaedzURfK9FFEQ6YPK4lXBUiU6INClDNVUqZ+f
SmdUn7nqTAFZtdN0KnLy1VJRGvqSFpmB7Q9EuHIN7VJBKlXr1WwCxSDj8uyDJaljqD7g4QUvN3Oo
qVr85qG9wkmJGbFEuqXmumKH6WijUrypvBDHDHogyetAcuRlkPDqz+q8c6EeVLL2NpOGLas5JXTJ
OxTVUZ3PcCkdnGxp0Fi5E3KqHumt9I8BS+MOjF3zE/tc62yVBtMFAgLxvMrVKmeSk9PSC0Krxz9b
Gn3nK2Z5jzH+Pfud4VAmnOB64tkbpl6fdk0XPP539wyoyJVkroGEFJyOleHodLsMKwrt6+NFsgHm
SpYhhxnJwWex/mI93QnEG7zzMKRY+AOXNyh0gqeoNBuEYN2/2mP6lxB+WLJVKoXEgGWOrOJ2mJ7h
Zf2gIiro7iPXql9ycYJ9MiCD+g2WSW87qxAU1+TFV0+e4DdYlMfOAVnpMh6oMZplbAQ66gwImQIo
7SgTA8AtoxvH/X5Ja33aMx9y5IyoCpTKILUotDHTd3FEFPt8nde0hsVoTVOj/gCYNraL6qzHVS7p
yGlljZHR4YT0jJfS35bNysaZ238hc3JjjAGNMOnw5dKJGXhdQDzw3SgMf1cH1quyqxtPQECTL6lm
cMlIkygiTUcCOMAiGnvBb2TrmhFY+cztWzLOlk3tkRJvbDVQO003pyKq6JD87FtSignpxADhrItv
qDzmpdwrQdKmfyAfuabD7YbrdOkoDkHgq/hN9G5TvIPNIkPcNQrWuSC0rn4j2tv0XDCC9XBoMSxl
9/DdPj4/t5bvJ1iV6ZgMA3dAr//R5kNGCaLTUTkys+67shz4Xsj2GOCDeKsV0tbCQ4qiIwxP7uIH
wkSGp7sTsx5zWfZU5b2VQ+EaA2mJ/tZfYqYLzWrU6GAUK9hMyaYCeab4TzcYPD5jEdE63km81c6q
G//PdPb0sAjyIhK5kaH6D3gLv0ovkFDT2CBAg05aKjYx4BaHUWOFN5EHcskIrzoXJ//I1GUCH24D
YCcRQUfGNKCoXjpmh5Urn/mYeXW1XN/BQqgIuH1EAFv3Z57DGAbo3Du2az5GcVGaLvtz8n0aBj86
jF5w8IkE8IZB2ewby4TSsW1YdABau6i6kLI88iPRSv0A4vJmgBtKFInwgQQoWvkZcjWI9mprgqf/
HlBRTdU1kLwyyEgyhs9Kq8roFjva6Cvc1JXz+zEdu8PDOssqxSEflbf2k95jL3S+4qrwUJ7BMXMT
mw/vbk4Q+Afypw/njUY0MsTTSHY+YcYPUp2yupZSmuUEzj1cYrTCEokHC4uChcWZy0NGx7PMf4s/
+N2UUJ/yMX0F1zFPtPazQWX3ZQvIYb5iGsiIA2tLxs3VaMDiOAsxz63ltjGvLKdDK8Fl56bdAG+Z
Jp4Z0GVWx40udb3s81V4wYfEqaW3pyH2oo0o+X88p3dwKXMvBf3YNVcYZZV7zq198aE21Fk+cW5l
t4fzZjQCQc5kIbIKT2Tvi7kXzZfBTWXISG7/ez7urW8rvECSuVnwJscdQFIhhHJy5Q6E4IF8GuJe
IPfCAJkrYHlDNUqIHAdBg8GDnjc5xJFLrbi12t2Wa1g+Vr3sStLKKbi8P7LbA90DCd0oYtGVHntv
aGjrepG0vTaqXxnzBthx8Mdh+iOSmZIgLJZU1TPYyLayKZr6FQII91eMA0ImXSk5m5uEayuYT3iH
Q9nVQO3nHEfqoR7ddyNRhHj5dl6sAgwSOn+B5RSUQr4yuVzELQQ5YFV4Wcig406j+SLbscyARDR/
ub6cqXAEtcGOBtfo5hF8iV3MrWtTduG8uls26Nc/kAeS9DVTsmwLYiJaDacA+NF0jYsfZVGeHHPx
mEfA1IiHWTYFTwlqBixR0eSyenNf2C0ZjccLp2i/Cf2DWa5yt8dxy/pma58jvnXiANqBkCh7yxd8
+Rocz6VJ0src
`pragma protect end_protected
