// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:34 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R/zrF4pd9BzFKTCMKWGi3TO2EjFggIfSEoikvrPMwCwUUwjI0d3OVJPB8LtH/daZ
8YHfv5zsh4derYjKskIuqVCOfG4gpoSUTURPlnK1cMHWVGOCY2qzlBfN5J8ad6Oz
rlxgtxiaSIdOyV9BAkAvNhvj6admiy21XNAV8I55Lmw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9088)
jQH3RxYIWnhXwsK8AKOfbB3Llbi1LNTfLypn2Mk1AEUat/YDP7fnRqkm6Zly0GPK
RwpTAj/EOb0ys2apCnPrVXxPyEbGhDam16HF9awxdFjd9Wvp4DmEL3hBDvCQtkyM
2DJmxsdjNw7Oj2QocOCNkwEke2W9UjvZMpmbOrRiamXGi6Ixbn+DU+EL7jcFJlwF
vc+vD1wiKN/s8jeohQaCmp5OMv8Q99qOLlEODL4Z3hM8cGrrIiXaaFbHVEnzhAIm
rOKO3QDiWPWHesTJ1yIxWFxcue6KuJ94VJDhdP5ylmSnjtot0eYpI4CDNllRuHdI
Q4xALUr8LkBIyrmeFi8oLT/JwP0726dthOPNv6Y892DEPihR4jeXna/z4aA2OBwW
6jWPUgzDwg10Yjjyr1K6gHh6C0yGWlZ/FBgINNoyfcDLHY78NEwwL74J+5y025rK
Fmodqi5+rnVh33BPgWGhCaJ7uK+2gF4jMyn5rW997naPxha+Ir9AFHNlQ3/eYWjn
fCwLD4UZ2m7aPIZRX2NT9aJPn4zviLA1HTZcajs0WhxwRsGBRU7O4UwS5pEzOtY0
i2f1A2+pLQYzaw0AFy1KStkeIMh5gz3Qb3bIShR2LLGD2dIbAijWFI0h42MpFrOA
cH1yRzqqAybD4nbvk2sHgvoCfuVNwrbuzQLJOMbD5c16HHcFracbfbEJPVNmJuhX
dUJud31J87p9nsXhKK2izsDeBvM21KC/XRbhFnpkKxfklQvkUnPWZY9q2y0/HnfW
HcEl+sMSGexg5lYQBDr7qKxRaeg3CvrZSvwlOUjKwaVLFSOPdFVz1gKqufA4nZX5
sS/wzk1NkJ2XJCdYIh1sF4GDTSu/ARZM4r9610yGVYgnCcrqXy27vEbSXk2maHbG
NZbiYgB+QRwz5/19/iAmRMoXqiZNd7g1QPwJuBy9lAF37wIJq/yk97RWaYgy9TYd
wk8Vehy5L+l72swj6/fivon/PWeLRNSK50hkyh5fFTyd5FDuNAve+YAvtg5JQ3Mg
dDb1QIWc89x4vMvZzZEfUSCGjaBwV/5egHo8RiPXaSpbpNxAhee/kWDrOpyITjZG
CXYKo63Tzw9Oeh1gUTErlP+F9hhmWksLrrqchEfP7+ZiNeSC8qAkbskymwhxGXuO
FhCwxNazVBS8YxGF8I7h8URhydxdhH9S2DSWdD2lC/uiUENrIzu0FXOdcEJmzOJo
CT28bExsyLLfL/1L+CWY4MGw7nIY/01Ns8jv/n13ts62ldT0lt69MK2+B8cpb5QT
VRxB/aDV0Ah2hPXiAUQWupKPZ173TGIXfGsyLqzlUFbkg7B4pM3+PgqGlLFj29rO
vcUCnSiRur4VUOZsBIhqrjtEj1y8GftYMCFa6qTMD7wOSdt7cZJjKFtS0yL8e0Xh
HWuZg1AeT8dzVXMwz3WYWVSM0LOgnLXwk492r6aaG3DcUvttBYYget5LgVhqmztB
/c9E6X9DEEENDKxHtmROJ98iXLmhZcwtr9zebn4VdiRoiUurQVvEZQXXxQpAgyuE
vfBfyxtO3gxjKJX8oYmYTBbomXOusjMBFgDPnlgs48usT92tlPcmKwsvm72yeU+m
NSewqwU01oTo35jeQk9Hr5l46jXjtFmNDoojRzsOr8jrz0HkHo6zOPq7YkLDY5dB
JlayUCiRYUg9sunJwFoqJPOLsk8XiUC8eyTtHAqBQzkICt2bFQF0Zpmeo5IHlEqB
6Atrf+j8n/9Cht3M+eHqxPdWdGMXtD05DL5CYqyZknli4M1qZW9Ox1ijLHGn5EAn
6Q9Sxm6izcfqApq856tXKSfCMeNOJleRtasaZwNxsrWslvJeaDCpF/Y19AbVEK2N
7Bdokzfohh01ABUj18yg1sYIM5K3vyvgbg3XGVcleo83WninO9YiDDHIxL1TpMI7
qxyMvRRQgkBgEu6M9GLRfY+68LD8pX+PBQRSkqKfSLfEZhWlraPf/b4FB8mI2L71
DsmSG2IQLg1u3Rufag85cRoBoAQRfVT1D9caXSX3aauPsGSinZYB22GJdklGiwgM
oCUvb0sHzxo6o+Zo4OyyjXYRd9oLkfpkUUXL+l2JkNaZDNJu09dPpaIk8TH2gUs4
qzyEmCraYZvfHZke6UwpgZ/jeJHwgdEL9DnWNjyypN8Nub5PEivn/EtDJ3pdPqIs
Z8DnBJab4UJ39wHbipzoG9f+9y5Vs2jqOfPN3QwsK3Kt7PJ4IzpruiO+Mkloxbd/
IwkP20TqFrDWeYefUgbMnCMeTv2uFE2XUjomlkMhM24QHVHxGdF9fgOhfgyZAaXo
oFvu9AI9g+OP4hU7dPC+EErREYC2nyqycdeCU+vTtudJYkq6/e+waz6dMwgfezWJ
/M+2tonQRkQFL9T2X2Xp5IqepyutBnkwnW+48U6NxBHVXB2GqbCIR9VIpVmMxn5F
SWN5q1zzBxm8UP47BhCJPwdivXviINJU3kDVgfAn9clviRV0zC9jLWUCQZPIuo+t
w6v0QzxVEWx7k8Ox72CebRBO2TZE7++LZph4Wj8TRe2XAfp2ztadKdSDVr/u8GOI
MuBjh4KeuPwI+EEHznyQQEglwJRcVtflowvREM1nr6dlLlngFcrXVA57Bh8ZGVXN
TinnMfTSJvnvEb2BEyXGIQlIqVSOt/uCPyUe/qFj1xklGQEbs8JzJVavRhf7Qdjz
kac/tBz9gS2qBU/73TctMej0RJ83nmL+dtxDwIM5GnxuFKEFms/r0bDNHzzQd2JI
v6bP+EV+cVx0xKCs8WO2pa5Me+2SlY/a4kr6dt2cTDjbdUeF1zLZpAhkkInI4f0+
WjD3pZpT0ZmjUPrnZNgOvLmfw2LBYRJes94/Lj2UpMvGpuQWBjxEXjnTCL8HSkH1
PwnIMOkl/LE27YQzOxYBFn3gTTn+ote2latZaDdP7SUKUyJOZzkvVrttuNECeUjn
Hy1JLI6KwiuYTH82FaSlHb/2T6XqsEwkAul8HDEHOObl7n2/FGqKWZtRR6b5z5Lf
N7pZvftae8TUfIOUeeUHS1OM6N3oA3jfVypIMyTOb/LNxtG3e+ApMV3jhEJzFKdG
iFewPmSvgEle8XXKSQ9USiW361UGdU45JnQ521iQmxQTB/Q0Mq5vGo0KlUmNLkbY
ntneCFido1emT4pymofPWweAFpV7osMPEVpe/NoRl08HqwZkKc2/0/oYASVl/N+H
t1CG2kyvaPcjydIM4OBmIWKXJsXF/uGrLNP2FB/FvktQzOqleK21hGTJA13cCCfa
XYD7vt0/pNjb5wBBxEiacCcz9RdfnGNzrffZ+lSvaxqpu9e95d2ylg9Z8uFAsMST
eQyZXD/dQ0MA3tV1vlSIkumT47Crnzf/pYyHGUQKsc9/66aOiQ2I6xJ3Y3XyGA4g
Z3BgjU424P7U1N0UcsOBGrXYANLWctgrWhUWyTHsDIvz21HGHoGi6fZz1ylJHx88
iwrw3Bmip7/h/I6auQAhbHSGDHpbNtgQp7PR2adnxzxfy7dA8Dmiw8C8b+aNojVW
05DIwwZvL/1BLz4eR7FxIXfNtDIT/keq7e0S2/U+DWZhHWEJjLLcDtM2fwupgu/6
nKkmKdBovpKA4kF65FB377espVaqiBkhhKY3FkPguCTx7ZrnEZlf4D3Z0s/hCTCR
n7ej2+lZuXMZAgHcUWtPGex7JLPKb6baqm3j+0yFYWKLt4TQfyT5jj0U8L/vjHF0
aPNZHvjVO3u/PM/hZfMaIMHcS69E/ZGGfEYM0lUL8kKmok4bU6UIKGzZu8Poe+OW
zhUqBup5JdQoesIx+d/epQV4Qk6/IDkpMhFtQivlw0az6nCFk5Nx4b2Y0xDW+5mx
dUeJlueqh/HnnCujLJyepMI8F0xpvXFBAis2NlELqPJCZTXHMoSw4wyXTXerwa0D
8FKCx1P4nQ8LGkqkUyxqoBdsmu6fAjm7TiVmP07CrjM3wvZ2aTAXrHkNFX+CKgFb
yjTg3tiQqh2HaLlvdjmiULT+RMVSiCpK6/J9r3e44rY8g+GG7jMDx6EooWX7yKiF
hH4SAf0OJD/rZMGaeeouow5CFNhzd/uyGSQiWfl12EVvEIHpNZThz88ruxfZiYxM
RYJHVvN7z323U/Wu5YBuzTa40mbbaRIGcTuxfa9VipPf3UXurGXIsqotoau40nFB
kpRSMpzz+qZK8yxq3L/MiKP6H6fEbH+K8XyBdDGDM0/uJGe5qP9IUcHdGseAJuve
7abAUE5m7TzvRRvOKTMfb2xkxLF9+xXfAeYQ0l9y3OSI600HnOmY/PAP75DMn5av
Mui9GYDEov3zEcvE599PJ3mMx/Oiqq1i0KQN/+LboYhcxhBpWqyCNazWP7nTRXIv
N0f/uZtoWbyH+NW8ZdaKxOT6TIKSfoK03KUwMJDXd8jHt/dauXzd/dtEPTNN3GRu
DyjTOAy3m7497jPGftcuNuNM7kSzXHRhYYuPlOPMZta2X+/0AzKm/QXbEH4nLZsX
oLUl4KrZO9Qdt/ZgkrKZ6GIycccMbklwiy8QEpj7Qp5C2MwxE+Zlnj/dVXFobwY6
YBTZ/KO7YjZJ5jE3eh7El79vEFD3C2J8rdY6mnji/FgO21W663fTvCuRbJuyYA9A
/prPtZrUZiAXfjwgnDoH+JOOSQQRM+wRaIAh+7kwNVQYAMCiaaawbLHFA9TDYpEn
PxP4e13Pmob9ObceqVCfqArxCl3b1lFhMe9A3pVf3joYDfaKaGvQVpcvepl7PUJz
mU9HqmSJPB6P205z5muMxZ4ia/dLRNpwEQqMZ6cmj4aDFVekILlzPJ32GRu1VQNq
DASABwn4/e5k5NH/BBI/Vt4j3Jm6nUtnxcSS7LMexCQOUGwIvn13ZbDTVbPMLABA
pOXzLYxWGQVb09SX5j2qGtzpbAdUc6H/pfy12qc9AdlPNsdv9ITRzStrjh1naC+2
7mboJqS5jUM4u1Iukxa9I/Y3/sd5ShIHkvOh0j3JDmc1P0m+/eaROKZ/a3RI3138
Ai0R32hllS1NHEI09b2W3FoX98oiBTKmJDmABMPwuEtiXTJKmkkc3Ue2qALdnPyU
SVGmdPbXimbwemu/cBgExX17Nz0sqCcjC00kUHgDHEHtmABIPjte4nI5YDZOfW+4
GQEU8PVq5zeLUOYFNFOxkOuOYdb6VViG1q5GgWcXqr4gJGffZshl1d1UwxKbkAMQ
mu4GWtntysaYlP4H2F6AwjaI3/n8bNRg5Xq/bV0kbMLPWl0RYx1A0Ymjok8kWsq3
yFjw1KwTrPv5tr1/+OdJhwQQgfnNcZpbOwXmoapLUwC8H7XjOl7nbEPkGE7oE70q
NyT7npsl7lKz0ILA3n64GUWGy3kgy0l8IwKhJpqpyuGmLRrKP8CjheRFmicoUR4Q
07e70sK9dm1iFx57SW/RIeloqaFu2Ses9So3iOeC9P32C97Ckt2gzWFY5yRm+FM4
pZrvFa/qyoSy6l3pGexU9XzYRy5g06yE/HZaL+7DvXTyrVpmAwyN2zHBBbUC8S02
78mHDe8fbh03BCSUPhfR74OLoy4FxG3yc5TFGP4PeOzm7sDPXy8hASdNFbbkId4z
fyUWSxwkZgkGReD5NthyXX0ALTwjnhUjinlU2jQptWAI+pW2NWgB9DPDHCdaBlCA
QI3EAzgItyzO6iLDKBYdo1/wRwHAqT4SzvVHjPGPGBlxpBs/005//2q8ynUwLONG
aRRqHiKc5UZZlzgOfZZ9EYI/noSFji8YnOEmOw77nwfZEdwg5J5Fi9QcIyIUqC9r
4tWY6UOpwdneIyc2s39MxLg+avoy+vDyjiBNW+obELuCmmckEzprocouDXR3ed2s
6M1qbAnxx5/2biCjDA0F8d/RR1B4yvsCJXniOOaL3xyS3yjopoSWzdWBocvHQeHr
u8YlKnYqVad1vKehLiKxi1s5nbYrLMc1smRXafJlfQK70bRidbD8L2M4o5mflqif
suU1+qIGQEVL9Eqe5iAuUud9oUK+nBnL9mRDsRTl1+bOn/pZ3g5WlS/nng9qcnoB
t9pfDhkhrd7Q5W8Q/lMu+tTS+UrswTwJaG+8CXIUMCLaXVlrFe9lPikgTK7fGuFe
ei48bmbwTEs0i0HJtxqEUN0BolQc5xvU2uuQxuuuTS+SfH6kuME66h1d+d/AFdjj
Y/qDWzAKw1bSY1PSt8L0wMnyjA9s7A5aYZivbQBTLizM3vfzo23QEAORg0kBRaOc
RuGKKPhAKVSbZmSlDyNxi1oyMWZ6VdNTrQIUPAobnm2xOQGjLXjUGIwlvAvfA8S2
SrVm9Vx7BLLsbTQOXUP5PKLqa1Tynkhrw/+VFYpi6gwLKkeVfffLQQNMy0K9xHrD
uJey1bBY3xN3BGkxzz69wdZl5bhssaLwnVFXV+lH5yphHQPuiBuNtcY44nNp5P5B
ZuKd9aRHYaBCyjnz8mdhL78YQgrP4NwGklErGzS9BtkQ0CIB4EyM8tsw/67tTzyi
Rf6T19+QMHT9QQmGyCDU73Zt2vGXuax/jN0yUvSEB97WZUWgBl3W5sxOH4aLvXT4
DjCltjXRjd4CKVlt2yvgHDJQaU64xyAjx9fAdOzaGI4jro4dGAyYDPYa+UMeH1pd
f4YOmQ/G9ao1iEAetF6QdH4e37ORblrSqRYAWfpo5OEC6Wd/qqq62eQhVLANgWeK
9veZQu6inujGRuqowj3BEAIqx5RC1kVEx1GEmlRah1zhS8kD9Yp7+ViRVdfoHnZH
i4LK6xN+6rZc2UfOy85viFKtFh6evW3aTj1fMEjCLmM34vsQlQ/s0AIORnFNEhzC
C3VonMDA/738AzftQR/3GNWtIh+EpCKPi+5K9usdIvJ9MGT1b7EHofNthkJlqoTF
XkMX6wES2mQVPvkXbfACE+pJmqruitDbKZbyEfPbHN3ZAxJs9SccbOeyqWhD0SGR
5lQwQ3HgtQUaa8/fyT7SVov+FVPA1wqcHPFr2ClRmPuxN0TXuxBnciOnNFvjWX7M
tB6v7p7hpaIfXgTkhlLJ+UAJSEokVwR47HvuG/eS4qcf5z0F1w1J2GyJnvl6Vl+t
cQARylTrIsT5WomA5MpryuEgVlflLmSa440qse9HUQ9Z6+qxxbDGKl406axGoZQu
40RYXjoG0lf3LYaoLALJQvCsgSxzm8A6qgteDLTBnwPfNy3QNYFwTuBDK1ZSeHrp
rTCpfgBAa31m6oVPzWRr226CBRBQW21DfxcV+YpALEM9EljJYNW6Uwg1jbITBPiB
Uxo6m+pYqut8qPfHiJdWQbcYIYPMnQHYT+IV19s8NOWe/N/pZnyaPBbqTg2cTN18
7Dgg2nz94nH16Hqr8Oua8RRg2wL1N65aGZWf8+QzzD3i03z8Eb++bypynU8qZxRj
2yCyr4WNLsxKL7vkdPP0CIS6DK/bCZTTMvje3Vs98ZII2YSpZ8xRMk0zn5yrqVM7
L5Cb+/09lsm822VsF5jj9GSx4tRCHVJxMilCVd9MKgSV6gS6213q5i4iFk2Hw0+E
4vV3nbnWiEC4xfG+WEq/oKbqTAqUmdH/7QxkyYvv6R2otk+B++de6FH/23fOLpw5
9Vmt8pEiWGVNtg721FmAcX8vRpHjseWaQFAdrCI2W+uMFvdhkdWByR7mtB3YG+3Y
5FjDprdmq+4ZUHMaxn/16fRhFCUaPNyxmu2w63S6ts+fpUIwky6da/hPE5k08XPM
nwRXuRKwrpwCH8MmkseptgCXOPMbemmrE7NmRftOoXVetElgOMHl4ibrVVJsqI75
9P3B57SnChHyki9OpgcsO6UdepS2abe88Dealff0ZS6bsxEJ/677QoIim9Lp/5Fq
trNv0GpyL2P+bmi21sR0vTLQJ6yKOBAQFU/TQXdJv6BA7n5gkNXOvbaCRRO2zwlY
HjLQ003azJE3HahIU+6KhoVUlBv/yD6DkpUCgb5lnnADDtIcwEiL1ecGdRu1Upwl
IaJLQhMtsNRI+tMmCCBKUQ9zSNF4nHfzoB9Klw86Bb4U6ggA6SBqfSQCHmKL4fjv
748wd/32nUHSpPU7FMM5b6J3y95EF/ELhUsPN9Jni0jFRVtHIUc4fPZ8z/pw6KoM
5RjQdGS4UbmPGoOSrzeFYw5Ig8gxEIkhmF6rggVvd6Fj6QsT4/lDJVl1jCee4dod
UxDqoBGz9Bc6GD6IllUx6FuRT+GDnkkg6/Duz5Tw2KRwlLl+oP+uqW4l1HD29gZ4
JQkb1pETWcOaYgi2ARdQXWa4BS5zyrE6/Z9hAI+n6C+OwiBX+wun//VxYJyJqgsU
uCXk1A3jMEQFKK6yZ6Xc7HIgZD80eidD/V/p3kWglO4HUF2RbHnfOPmEzYOq1vsn
4Ipr82iOGiwgLxPFweqP7rygPMYYEF7kD9RbZMhG7Xoimx4HruSiyjqdL3uwZ255
fKS9OhrXT0tN0SLexJWKVcW0btzx3MzZvt8np6tHzlYIYJ57h3ZZFbI3fTJyV894
fMW+IDvkAzfPEaRRdOiMeRzEh+7LJsVpfqpaJ1dxMIs+jbm+KA0YlF1i+AP41mtZ
i1OP5tXhBw5UyXvQlJ+fJXHJt0IDmELg9/+hY8vJKmHwDpsdZKrlb563Ark7NWH3
Jn6VUsuYwHzJWQKB/LpzwXM29Q4/uj7xyzacHEhrUcsjogDx5ZkiSzjAZYoHeguw
DGWBxuvo5Yjh2/2eCgYp8B3HxnD9CRzTJhSuJ5CNqZLXKFB9Q7jflRbWBPJk8T5l
lvaM+Yie2zUVQY5TiOGxoX8eFlby3vS+6SWWpoEX8LBsHRlNzxLtJ8P5XzYnxycZ
1EOYAMyqCsfyI9W7qDNtFhCFCXgHSpnVCMSkJSV0zpM6A84eIkhkt5R2KwaDij7Y
+P7ghO2h9kRoHP+N5TL+sjsjOMpz4SKO9zdASWxRs9kFNcKF1MUZxz/oIMRKlS6w
+649YkeiVvjS2zm4AXJgYftTsmfU2XT+OhQXRnawmQLFwKbAk+dFLLXO6NHNVweQ
Tn3yDgPTiUz5OrOyVdPcTejPX5pAhiCkBy513382+HSXsLOANDmCYjwmQvODAPsF
eMhRfiReX5YLdZrorkCJ2ovBwTmoxQZs1WijnTzo8vYZg/vPIaNdNKXCvHDqlV2n
8AjnE7bON4vFc4Na6lROlm6vwvc6JEK403zu51gzO4bdU9lQQiXN9cntiiyxHl2l
fWZ0K+7qUAcBkjZZgvwXMrH8bxS7p0nWYPTcHyfA699h/ZQxSWTjBIKYAKOzqXFE
O2WS7cg1SGKQiQGioLzkvEwc82VPodktwpOZJhJwE6efLyEFU+Egb4g0Cav0Vy2Y
HcyntTrheVesLRYmoTa9I4OG6WmXICouITSSNuTXrvFCplS0Gx0HMwrNHBV+9ZvK
EaOkIw6OznFTapvwTXADl+0KrVerSyGvjDCxFSfbTPAwAf3jxAUJoY7C52+1DSUw
+uB8mOCbO+JiADe3smdxKXbSRWYbCaSb7Vz/e2bZRUimvLFKgQ7kJmmo4Ll24IIQ
Bjm8owJ6sQqwCmIGdugZrSrEYAMGHMvZu7p6Ab1uiMOKwoDEn2D395+h13fL13uQ
HrtKovESS9ZaqUOJ4iLfQecqkR+NqO1025OU99PT964g5kcr9RNdZw5QNtWxZdvV
U7egDhRIwGxleYt1J0Xlr7a1DCrCoMijeRvE7FjIUbF2CFinouPH9Wl1jTA0Qnwx
ZkQim0zjncD043l8+sXcRrd2rdY3gkFlsaLVk+QbniQ9Bys7Lllo3GFnyqgELLip
l9ZHe8gS35XX+2Vajv780qVEmZJsSTputFK8qefTpyc2rsYaOd+tYzZ9hWoRVW9k
TIP+f9C0wubpg5dpH5AZzTnPoVpQIGxLCU03Dg9Bc1wPIL7b2pjtg2ONvCIZcwsV
fB5aC4KlZSMa/sKJsvV52andVb9M6GKlm9T+M1Cn0GWzBkAOLxOkQKCks1cSMpsg
nfEDtC+ZmdyRUBJA7f6S23z/cQAkEbc+dH90yLpCChBJsA7NC/IOuP5Pk4Z25kBU
FKx/TxNRdl+brxyFhMOvCfyYleMxmC1RvkXBgI50Z2p7I1AVlUvuOF+2XcDAACfu
A9NXZf/KOPeF0OD25t6ofCEEoWP+b8wW/kRMnfW7m25+S6z3NKHEI1QAL3c7MEix
Ktwfd7oKUJyMKlAOiMFArtInXXlARxDaZ/zbPtjAmp2Emjpu2y8uYTBBWvJsBbdS
kuAkQgyXMbgu7RuTGoFwDE2aLi5yE04br/B4+TJxqj6XtsubSOkRQhMBlK4sQJKm
I1MSaytd/S6/Sin0KQ5J+FBk/BdTnRmE5YD/9cQOdrPquslN3RIMpc2ksHMadiV8
vDP+7GgCe+0yAPLsb2ECuAfmD5PXEo3PqRBUYyiCdd9NLeLDUKCL6ku7QsLcz+fR
Trmg1TFbWWdoD2N9TEmWTaGjzjGg11+8XJ74aXcntnn8TK1L6YlckBLALRMmUPIb
NwJ90ET+2KfF2TBnlKKmMC6I0q0vXQSqDkK3IADdQ0H83+WC3Q3hu05NCnvz5y3D
B9r5zOFn1vPDihKQjwbMubVWUX9cRSeN7PUwXsN9KiyZjjN6jCsi0t9P+4WzMaV+
U0h2+qsEog73PHfLVbVY029lzjehE27XZCwrfeOVP2hfqsHthFFXFgkURLtyHAIY
3+XEBulsfov7ul+fPz88vIUwSTTAJADRpNrlz/raLCyMSta59kWQRxFXdixdHzGF
TnFi4T5tYNw0RyRoRDab4Nv9C3HWBfc3RCu5agTeONDLa5Ylar35BLaXzTwYFpvh
Qej9L89YGm6cMDyc+VrEw0waHkXp1NdFitj7YYNgg3fJcjKyTfakc6VjV745uVuR
t20HoAURqsxfZniT3W2jjmSCUcUAP17SvvVD4UrRr9hL7qFz11FPCfpQeg4vmWqK
MYUhHT2yI+tjoJJqBUUzGEZo7JlEaj/uPbooIJAQguqkEF/nBtOGGpsh+FC08Y4X
q4Un6zq7RIm/WTZy0feQnnwEnKrhJ1tZg+bY19uasq8MsMg/JVPJihjs096JdS1T
RyT/5gHbiPsDHijpyvj9ryHqWKsZ2l3/h+edqFoGoDQBW9jesHu8vhH+ZY95f5es
/idaH5HPM2+4HcD8X94SYWqJI2sV0lgVZrUFv2Ge2MO+g4pqSB4bQd1zZQk2Jjos
5kpnrLr2mmIJPVtpgFSGd08wTDbJt1J0TNOUlss8Mhlx0e4Vp8m/pZB18Oz3m7KM
gElh1CsdxFHJ3nFLJh/wbIUCULHZwRGvQCSNRRdrZJwoapB+A4ZEUBr+khDQy55p
WWUlNTIIMzZ77MfQZaGEkQP4NoWzJHtrso7HUyMyGIqp2cXELXJpjS4Qbu0pWgSO
DFidQwxoxtpYUL7O8CASWjLaeRs2znGrra1TdWGEyfy2Y1Tn7N5+y8A2mujTwALe
FfGr57OgzFNOG4xseN72gw1bxeaJ9ChTUS+Q1I39tLJM4bQ8q3AkkLdjbYU4LLGD
AcB7yTQOltvJFDD4jzQLgRO+FRQBPSTRSx/F3RGClof7kXNlVBQwrbVpN3+Mfj6R
6Z1shHduqiUFejcNRu2wWKIeCpBwKQLMK2FYBqpEW4hDpVz9f7otR6CvLiyhYUGz
NZm4qkW+SfyRZZ+o7j/S47jFcZnpkLXLyYsfLBUMiyjxiXU3pEp3qZIZCpI0kPX6
EBWCihtMGm9jIDnrjP0YIQBl1n5vkWhPh73RA9tdOtu4pAwpLR8eCyI+fHNSNsiO
LKhpCnkUKX0z9GQoGvYazwWS3GMSMoYZd/hXf3OGEmDTZ8LEi1mNbTbuRhgroNTh
LjvjcRuDn0SJVWSFEK13wG8yTj4BaUl9XwF07G84T7XactkqCGmDzD8FFOkn4xFP
SgEymQH1nhIRDFF8l8OZNtuXSv3kBoNPfVbkOkDOPUsZdesC/YikI/ZoXgjYcSDM
NYq6vPkvgG7dNOG6hva6E4dpEMFYosGtaP3jMV/5QyG5Q5vi4K3Goh4vbUQlxC0T
crtVf5T+uQWknTuWOTn2rKxmwyQ5v7dwpL9dIz+AN15AN50Vidj2+iQ+5UTS8MnQ
QSEqGkSdpe475TKcWfP6+T2G1FKBTNTdxipjWshowG3vUUSxVJC32cN61tf6G/9F
dFl8N3VoRGbAK4Nenq9+pg==
`pragma protect end_protected
