// unsaved.v

// Generated using ACDS version 20.1 711

`timescale 1 ps / 1 ps
module unsaved (
		input  wire  clk_clk,         //     clk.clk
		input  wire  clk_0_clk,       //   clk_0.clk
		input  wire  reset_reset_n,   //   reset.reset_n
		input  wire  reset_0_reset_n  // reset_0.reset_n
	);

endmodule
