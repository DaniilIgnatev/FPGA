// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:30 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Y39QAObkkm2iWmSFVHalwW5YErSh8tzmPmitALotUNAEBFdPJcif48Ml2oYRw9a9
KE61QaCiPzeGicptYR2xPDrIxHYPPpKs5dEs0Ihvq87XWfLnWeIyxyBf/5Vk+Exv
dZf42orSGPdKSiIxXPr8iWlHzitDU/CFJLcqGpN0z/o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 24512)
5PTF0qs6CURO7QviZtaIi71tD5cZSz2xxvHUV85ulptOejzgxnpL+mmNP2A84bqp
sFn6KRAElt4/1zwIwcRgqIfTptBD7yXuxTNRP9VDsFY1LpXa5GEXP/jifUD+LbD+
OeRg+m2FQo1gQltSk2RzvA+7H8vJVAhdTGBmAxyUCPMFjULlqIsTHkXIBTRQtEuT
rYI/7I1tk/E81mejz+JFXrUVY5b+gVrWZiNw7y/UUdJEEIuXDXAr2dewTbIbyYKN
02ruvs+KMRRCAHmJMn0hYc8GGq7UMCOsg9PmC9AMe9kX6e50riPoqwcHatW9sKHE
6AkNO3U92dKOEVNy+kGdsFAwbO0dFMVV5Opl0MgVHmnovwOuZz3EOoH/sMFsFEt1
2Ae/uY+4WRCDwGRyqgHIQtZSpQU40G2ux1Qk6WMaEppF3QxpIzShEIfYf0H8rDE4
N4J5vC56Rjr84gxvK1bPeU/5pTQwVsKVpudFyOQ8f8PO1l5tSsDTAM093YT1/bOj
OhMhmdkySTRGBwm5FDEJvYVN6KeQMR5i6/W6XI2hCWQqZwcWkSCAV/zE3WOEu5Ta
AlmgmFHFoQza6Wm2djDNBCNI/8Vi2ns4SsH+A1PdYH25mnNO9r95VIzlLkbDvJYQ
cVkMRDPVAdNQFjkE1skmY89QkNRDzD8SiCRsHmswqwcj5eo/TcPizk1mty0xwnhd
T3VL5ECgFQeOlIAylib7GjR0XLG/3h3kweeCI4yi25mVumBhBA2RwjwOFgZl0TAA
pZVs3FNK5Lhq3Pc0ii05d6WmP/WsPomcytBrEAiEAG9uJMGPdqcbMptNFWq6S0Ca
6ZSsqk5R893eNprlCOysMvd3sm0il8VivacYK+GNzE2HnFI/bsTJKB+mGNVVaz2c
n9KlgfF9zSktnlJShH5k+2ur0/T9AmIXuXKgrngPyVUSQXVthH5+WIKr0YJwSeM3
GGRAzaxSBtakK6zWztn+mMUigv4fnKNhrhxviZ4Qej2si5fO2zOV1WQycIsyjc6g
Ie3BnkOhLgVMyoA6T+eGVN8oGW7CZRWfm9yldeREvXoO+D+lkxQChO7tyTs3w280
eNSD5B+bk0U8e/BBvAoyV1wLNPhqHZhSdXMqkfnmPH2tEojj8jI2//95alIOFXhc
VBTFjyrQ0XM9qFNBFRxziSVX1Unur69bg4Oqlgw/f0mHx3KMoyAv14UIQRwvZVbx
mbekKgWQkV2Hkm40P5NyFourlGA/Bqo00XuR7r1CFCHzn0ydqTGSbAsiBO8KQg9y
DKjnRhJL4uey6FWyI0u/SEcgUSILVAOw4k7Sf+nDJ+V3JzH2EViFS6gu2uXiZDrj
f+X0HvNLIoqydjSb7oQvfibrkB+Pqn5ssRJK7ht9PGAVrnXND6bM8ShSPHyAOjOt
oTcWgimhaollW+dF/amQgxI++iV3LOcNugXacnpW4s9kJd0RJDbEx6iEbUwfuC4L
w4CF5VJ86LJX/slTmf27udrdcKVBbufAiZDVB81dkpgNPjpzkjiX7PF+bhgXDda8
t0JDjagrI5TT0BpGLCmGbpeI2pu/wx3HpYT2KxaJWvuyyA0fGXpsMSr2IV7tWokS
whk1PG2kksBiyRMAs3ZymiOnC0zZ67H2By8s/YlLN9GqoKy8+ZqwR/VCOMKat97L
xBcGbuBnsoThGz/u265VyPhvATfGiMwn83OvM6Jrq8C3rDZgv4nRDPx6V4qyjIdg
htjPoGiMaPcemKWVt7tvGkb1zEYJPwqAeuSdcx+I/t2mpodR9Rc9umAVLGRtT9vx
2x380xkOwd2sWscaMGvKDrqeuMxQLiwdWd3bPxYhmTQ0iiwWcwvZYja0DpCY9LXV
IVOhX/EopB3OoQHub29qfDMr3Wr2qo7cCA1yc942kXVtzes/mL5eMsxFhWdgDI9S
O2+M858hxXkBpqcm1fS6H8AILaww+ELskmJ8V8vEigBmQIfHg0lE0hLdrQCA38zY
aL69AJZbZJUnQ1I5Lz8NBLOCdackoFaMvtI4Pc3uDZ0zhwns3BvwLTXJmFCDQzdN
CgrNxNuAXvi9Nqx2fNI7dfv2ECDmCSxxVsxvkXl4/CqlfqUvWxJbzBOGG7CN43+4
VMXAUKnnedx4hYqSlsgZGjp2Nxpz+TytSUYxQW9kcqkChinssFJg0041rEX6hVGi
WmkkwnGEkvWpkt1lVMU0PWQqrrGEOKfbvZuTNDLafPI3KeXGDZFbmcTCir/sP6Of
3mWa3rHKNpuORSGHkkxyoLRiygPZ82kYBtwiM+IzWtgO7s1UsXsVC7KPHzP/sK2q
cIbr7quAT+hisBmEXlCWHagOVXoIBlvynu1CgoQjo2Ya/fGvCUlCePjTKm4Nsdha
wLJq38qb/FtKqK9athyOHyDeo3fRdXWhPpswKrGORGx3X/lQFPGh+0J35F5rlse3
sixxfhhN5IG3A1eVjTckksBU6JQoVCX77pr8/hXAF9WZNRoND5waMGgx1J4HEp56
9tEmwtbQchkti9wqtRdwp/NyraMo3Fcb+jgDZ3p3S/YVZRWhG53NSDqEtHKEsDwg
SloYYT+LHHwlMZ7ZL+70AgJQCV4GD6DN/G99MkuoYd2aKgS3mogsSTKzJVJ7zPCt
ndQfDmyydJpeYu2K+dcEVXWowLMBmP7OnNBpbdxIzOanmJnQFX8mu7KoqcAUS5fW
wafzhlr3aUlFqe3RTakBn1U5FOhrErGL4viIDwg8g4+LWNHFLoZ8yizrvL6KABfw
R3j1hRoQ3d27aJHznesSun2Gl2R6MpYJByM+HHPkIjUXk2Eyz2r+2B1QDlP/1eeZ
6siv16Zns4nyzWpjxRzQ1pzHb2spIxE2U+jSkjLEEwoYjeGGhVwoqoqQAkfR/AIi
rRpd+yQQBDMTGW32lQakpf2nyCZwk8XOssyTdDI+gdC7ZoCJZs/2q0tizKYXEowO
OQ62R/9qLplGtDeCSVdFF7AGITw9KSXPAXffaK+xM+DD249MQfHhib38eqDhBVSj
elyvqKSnDswkRDwzG8rYHVIUfh6SK3AxL70WYxyUqYYy2wdw1iado8Pd2Z6a8sl/
1lXc6P6C9nrfSVPPYm9LaVwHzzoVlG7JQp/bb+veBNZZAn7hCTZcSHxBlVLUCqZ0
IQ6LV65eQyk+zZV2/9n10l/x7R46s6O7hKFh9Xpndy7vJ+I9KB9WKv3Ni9S2Q904
3biZQPQbfvhR8JMBlEvYGFmNrTx/xt04Fp9EzUz/5dLhLVRSBQrZQ+OrUvd0AHnJ
CmQWoLGHE0MjRbW01jPOd3NLzUSsHvNM/yujYRcScuezCglF2Blq1uYsgJtWr2Di
e5U99NEUIq/LR5i6uN6nhmaLBbC4tn56XnnjeZpK6MOtSO8LQ6kSejAOK9FLjL9z
RXYReM6YOe4+aihAVLePdguipjkQobtYGWtQCHNeAg89BJ1G5ApjfAIzkXYbasyz
2DeU33UBF4STP765Kh5D/l5PE7ThA8wNNIPF/e2P7hU7NGBj8r3F5waFJWN8910G
HcUgWCzs618e2+wD8ezDg9XhfeJcPnHlMctca0+hvsjOpCbnsAlDmU/8pS+gLeLd
3o/lhnKfT9aPORUpthxknZyOfUfH9F0tBmoldkZKXdpk8cJDMttFLtbQxCpxROQC
5AVfbGaxw+2oT6aVlU4MLUxQ8DsjZUB7EdFriIqCW/cygedn6G7rUxGDSrgKg7SQ
nseB37KwnqVR+GwH8otvPeTr4ZCYaQPegjIM+qjK/nVOsfdee828bLReRtW3zaQ0
z9BroykMWVJKzYUAN5JoKF2qMRhhx18C/6RgI0E57Krmd2Tdh7clWGpf/HT204of
1QAj0oiqv6G9kXowE/FbI5Z8Xi/JFafx2gPJmmsvIeN3Nnr1+pCCKzUU7NUqxtbO
fisUApBQVx9E7kMHKI6LoqlVnJJ/2jDcPz2gtlhVFGTPDZhd0wCb05NNLS891SL8
GeFISI7GBsKJPRtRiAFVRxwMJkOYLHDfaZiZ0Sfq6aHb4TNqBVVmo2t5dMjEdptY
mtt2YvYiT10AYlbjV2KQTMzpG+Umsih5PwSLGeysZvTml0/CC0x8xpQo/k4AozcY
IkgSmE7cKS0Ng+cHrLh00WDqJBlZmfs5CVOURMVHGcaTrLzIUW/MO/4lUByEUZR/
DEigVfNoPW4Vgc8MDdlSuUBvw975MLRT/sifLL4GyqTjKaWAShARpA7fE/a8Se43
/fId6HC1qQ7gkV6L5VIwrddK0BHbSfshM3V6zJ4DBjqczBm+MdDHi8hZQlLvpzr0
AeCeqDQynvjU9lsGJKaCAdBeHbZlDhTIZTjgsEHSnswZ9EFxhe7xjQa0qAlgnS8Z
pFsKdfNZSsLUOcj3Vc8cMbp0Si0PGOnEp+JrVAezwtaXNHEpNaK9edRpqZZpUU3p
KzNcq/WktBseFVWRGPI7DUDIMWfZpI/cFV4woGreLL61lVEoK/PAC03scl77JjmM
nqdQ90ngYzia/dptLxNUuFgQEu2K5hjiPN/f+1Ky0+Iysk/YwA/8urh1DnWNdb7C
kZtrTM5deHsCMu4gmaWMvnfsuDwJAWSyUe98gCdxo/n4zEqPPnBqrgfz6pCj24Ng
4B+TILCYK46gRhJCeK5B58V4RNzGPoxW+SpNhoZurzoSyEuT1mMIzIH0i5RYraPl
gKmsdjsTsn+Y+7/b0FV/0OGqcS2+1mCKoZVdShadYtzWdmSx0rkCoeM4DQAH463g
Ky7VhrytK+q6YT2Hzmo9wf6gSjOSlxdCY8m9edf3cVYqiTpIkmYI0lxCMLQR9rcX
gF2fFqaeYtDmzPdzasPDkAYevC0Vzg3JRGGxl+1CMOZ30yxph3xiEE6niSqOhqSo
JqvAZtbNCJjfLkT49stPVPJUobk7hW51/0tFw9Zkv7F/Vj1ivrCL/cb6GEIZgdIy
sJxpdshfAf7QjhKzx5dRU3wGoQz/fCvUqJAyBENSKggAazJa/7zE0cIEfrbetaWk
ELaROyIuL4PurB6r5HasKG/7Pi/moXZhg36+Tvd8Wl2yHLY1r3zmWiqcHH6/MWga
CIa67RXs5RWAz3fcj5CVnUHrhKda2cGl+JAF2JK87GyfJs8mstDgYDVsO/FxvlPE
g5BYM9AIC4iKp/0Oqxx+gxAUX3zGV1qI136jAP0CmzK0O9+HM1Bgx07B6dU6DUTT
eJ1TX2W0yF204ipmHVmF+wzUmQJV5VsVjBe9EUIoGpxAC6yu+iuVN+L6VnrkmgVv
mIsXAZ2p7548sOdlJNM/uiteu9gA3g8379sU5vL1YHY2PdlOb8+gXwOKlI5ST2AA
fxGgG5MMMFAFsQ4oFwCf0kheiTayF/POJjq7H/dyF7CVI7feblOdutOpEJe7gGhr
pw0vEpELHFoJAA5FJxOD2TIDC1p43dZvvNb1+MVNjoYN3Fr63uZZum31CGICTErQ
qTuFy4a8aYJwmvy+PVXtX/WeXivpCrklMd1CBEwR6LuMCKidTXdWln4ZacR5B0mO
Pvpq5LIhL36fT1E0MReAnth81BTydeYMk/SbZNknlBwtjPg50PgdS7Hvp1Z+66JD
QzrpBg8V1e2U6/ynz16KnB9f9SE7y5Ky12T17bDze2ItD9L3jeEWr4L2Jky+YfAn
9mF364DPDZNPRZU+Y6AB1Es0NzdNu5B+slcrmjAMEpCZxhs+nLd3T/A5ZE3Si+Zd
TPpn8g4Rff+fG1hHkZdsfU70mm+Lr3N2QgDS6ee6aLgaj28HWSF975IYSKHYd/9v
SbzA+108cZlA5nS9vqrzUFdCNQWbuVmAkpEKDs/Qe0RJ94vv4Lfgr009CKcc/D1/
nw8nSYgCoYGWHT52CAIV3zio/lO9t6PUEcKk9mAebd1uK3j8DaDkqXXolx7oGtvl
y2WsSzAfIkmbxmqx6RrOJgq+58BDan7lSW3tR6Jp1lTFqyh97OYh3Q0QhYsUGNuT
jHkhlHizO6sy6TtLfdsEK2YaX4tklFB+J23iotrukY9Z1ncgceZ0A89IdJROxelg
K1kV2Q31zKzVvapPWz58jJVMowE8YIebF7bbCK6L3XRsSmowLfjdhRDO+E6P6But
m9R9WGJVKLCgO3oxLbZO2uGQQnIPO17vx/+E6DKRVz9ouiadqdc1iZvJTg7oqTz9
Djstu37RQ9a3s9QQSRU4X1mMLgpQynhnbYKtWgRRb9fHXLnaE8zVZqIq7DUVeQSB
B/m+lnEyvbeUGFjxuXTSe0AyuAQ9Ro3mC2J7wkP1Nhy7T75KXXjAmWlz8w7bluos
FfNTvcqndZZfBWFJ+hNu2Zcz5diGuAbLxVlnEyuOcJ2oMlcFe5KRQkAmRD6Ozafx
pUCQo8FowO96QyNYEs6ZbbfdYXKm58ozHsLvR7IXebpv0M/VE00fpVRl2Gn5I+9l
plOxjTNU4JsMWhTt2WpQl+hZQgopm6520u3CR8DH5HCohWU1cojqrlJtYBzaDX1J
dWwVU3UW5/vtJONT6d4sLncxgUlF3T1a6ZCk67ebz37QXqY7rM0510nPLw1NZfqN
4haGgqJ1haB3DdDF1ktAjzyuIMrkn56j08QhIFXwPCdskLvbXERWsFdi4fodsRbl
uD4EjBcnHlGk9ihGww2m6ugv+CMvTCoenqa3LJLjIq3UY0DABbZAiSdg40ZSeDpl
+esa8NZ+y4Aq0YXewyhGPv25MoDjVH7MgaOb+YqV8h8584f0ysRt3JdEKpQIZnvs
veP03Z4gn678NH4+1nyTVQ6PMwJeMSGLqWFQyXooMZxUHQWgHVfSkNsBmFQdtcBW
m1espzpZTY2e9Gc941OObgReFHVVuoxNWy9bAKZRgpBRhjHelavT92eYDKUaIWKS
qRj/aTNkurMcx5pSLHdFkJgeYY1aocd8+VHRhUWsIRYtQZG9qn4Zky7BiZsgvK3J
Vgh3VRJffULIpJCzoHLIG+vfGjlg6xfFXi2kHOVMA4J7juBEl8W0rfwGQeCCPtxR
u+E/TGssr9O2BCpTQtEo11xAbDuxj+IA6yLiAi18T7D2HGt2X2FCIkMZTtpemM3n
xqAj7ZwUjIN/Qt5tsRFy6SKkP8sM0wjUKfHsUZoGTOCxIHFfgYj4K4rGvnFfAlgn
06lfSJ+Q4qiPxVIvY1GMLzpb57D1iCsXNkCPp1XpAeaQISbCP6scr5ncXvFME+cj
pLBMTk4DyPt5L2P9CydKpz2K2UAnuxePYNwfrcwobjwFWSbvCTZIlmeSdZXdhJ7x
kIOjnVJaGo4Iukj1llIiruGJneG6fx3dX9FW6ek2trYhIcVAg2DO/NARiTsocq1Q
zIzM+7vIkozT0/+GaCnCnBWFMauIpDVQG++Un2eH4Tgv1OiNERXmJa09pdxzEylJ
n7RBNDwvEjPcetcVlIQI2naGVZlZgP8N4Gacd7jGjn+F04mR/k71AVbUr7iX02Sz
zL957Y+iXxh2ovBAl+sUcSM5MVAKUdtcWjNXQYBrzrDGRjFqKX/QtywUJf40yHiV
6EI1N8YAoVbgp40rrckRLXq2zQcCdWUzjJcTH7Jr6M7oEPEZ8yT6m5aBZKLHpZH7
qwTvCDVANtYy99QthuR0PGtisCrlK1im+5A2W1/d/SC6NUiCLv6XlPZ9YRivkeEB
gQxCffSLU6KPt3gWljFaKvCpBVzuPzzvZB9Ww+2bXKXWET4ndzdXAzwEz7TxsATl
gWPj2RYAeO2LNZNys/LO5AKQ30YBFClqeJZtNqgy4oVQhxlozFqXtrJWpGTzhnaN
vmimzJzbExOvLoY/rkL0x29p/Pija/nbcEm3PD4LMYrcjGdpd5oo2xAM1RqsqNnu
1gMolrRzqLupPTMoBcdoqNgyt/8+3C8eyF2KI4vuejFP5Vw/LTEj4yRZBQCeepGN
KZ/9aUV/KJdEbKOu5x3ALB3cy1TPanLvLmu/n7DQ+fOJAK4xLcyFL1en8x5nrzTY
tx4fF2ZZRHzCnVmTaLICV01wP9jh8sw9IpZImz+BESPcGNxsMOYOfB5oXG1T1xM+
upafnIZStcuJpGUlftv6dgqsHuo5HrmLs+oG2Wx2ccTJLjpex5GugsNPVBpZZiqT
nZjCGrhqMDOPMgGkIefCU9kt/2VhlKwCUf+XqOs0gCxQCm2YDfaMDh03dnZy++s6
iIQ4nVlbtvdHiXv6G017FXM7Q4t0bcRR1KAB/Vq9kqoDNBtSlIGHnPQ/NlPfdiYI
fiQm8X87KCBwGhSrPmpFW6+XKAkDLRJ7j2pIyWMX8r9vMnTwzH6iMloHUU8MCzSj
ZVZfkEMcnofG1Ma8NdHtGVcnagP50fdg59EnHADfOD9r6RLBA+LzgRHMeFdqBb0c
LjBPnJRSlDuunSHpj/yH+gHbfOvQQPJGIwYz3J/3JdQGk3QrDh4ShSqsESmkn7hC
H6cyc/qR9kdcVv4Y9Ysv7IA0aIlAXQ2CsSwscAzOpfwapcYiuldjA8EOrzpF0c2T
gwL9QpPjs3CEcQ2RWWVmbwP2j/5PGZ0zunQmSBmwphQiAKWsLiMaKT2E0ByApROn
LmMN4MdFK3WqB9gGeJNqWcn3qjaKOonN76A1SX6i7U6zPqLHvCKUlmKknxA7pBp1
h3bnB9v/4lunhLZBfd7E9JNJsx4vNQlWm3w/PLGtY+P5Yz/az/nv+lS1Vdq6aeE+
NUFRjJZsdf/xK9YJG3iCxD5BETXxNh/1J4Lro46JEh3AtR4RVzHQtfTnrmqOtOZJ
HqCnlhOtMNWWqM7vL3QMlnuM9sb1OkIEA13o8qUpNZtOu+qFumMEAZJMEC1JlF0z
30TkKCbKRfcbv/gHq+Cb3SQe/hOfpEH24xa76NrQ+Vm0Z/nKyVBNJSOn7yVNxoAj
ljMV32qgjqrJrkEmURFj9lhNrke1jyCICde992ihD8zLSg7fLOcRZJt/UXkIbcle
ijd7cfmIJ7uzlUXr/mym9hDcAaU/pnQ23MV27Ho39sBTxRfYsH1gBzUmm8s2ep5U
yOWsZUeausCOH4Q0gCjCwoD8nu/judlBBgoDInaLVNmauYIqC2Q2eKVTShnWUa2e
FpPMn4or1FIBUio18NaMUfYgtv9JV+sLweuGyGmqHf+YenpzmHPbTo6+wyiCkuRO
ZPTH+IjUJZzNUwiKSYYI9Wr9CPjn4cXVwtY0xxACUPEaGyMjdnjl+1KVWFew3sSs
/gypxZ1M3ViIAUmUaJR8v/mVVCDODabWvH/dFDWYXAWO2zDmsgXHUgmyKQO5b2DG
VEPzF1AwQC7SVlzpT9KAjA+QMvk6Ky2qPsURxHxVM/l9J9vOr8gX6jS3uTs5FBp/
Ai9zaIGY1moGyRv3rg4KMg/jiadeseb53DERLXrd2l/sq5PVyX5PHDWZHcj/34/D
iOKKNhe1Nom2Nifh708W6S69U5qwzSubEuX3/XQAqE9UJhxWBN36TJA9PMWsYlVO
5vxBHrd9pwgslQNwgmCqALBSvc6qCzjiRfjERQvS33QhxOmc6ZRqSU80LeBqKL+n
vfyzD4L77UNwDEVBg8mYBNJODR/+ySvvRmm1TJU3UUbkKFOq+aiT6sMQER5+fciX
VOC9lcrZ1JcQjV8zvh1IHAD3hZBfndGaWNkkQPjwDv3nzzylYug6ee9MimiXNPBW
JAPYHR5+/eNi32a5JAtDCN4hzepXzCx9VdIwyQmp+xswmtOxlqfZaiG45v8WZKRs
gbCnjHsUMsiO2DkC1W1kblHZipPwcB+Jdjtp74UYDx+DJQ5c6r8jL+YqdaSPZN4X
ZMQRN4AD/P/KsJEc3P4bqox9I+/izMDmn35Ca4ZH5j+C4GZg+8XmG0MXQWihri5B
XQYmcR3kQplAKMxOOKxozilvduPB0iF9DJXh2DHzwt31/RaEdJWPoSZDDL76FQ26
0pYcoH6Dr2Vtg2adR/LyDCLGNTEJV8dnGT54csMuVI2WvE5LsxQr/T7M2oSXxPaf
/3PMmzyWztJYb5/8rktpPQ2EWfNswPCFK9p02861QqcFv91on7wSTbv7BKsi/W9m
dkp+IjMJT+kLFJoGZ+4TF5ZlNTt78NCD3XlGIMCMAldGfWSDukqbgDHStABqBFvt
Gbqfmq2MYTIm9GmSZvzZ+6m0I499MFrxN0SCjF2UVMPARu2VKhZ6xlIWGeM+TiBu
Z++13OYPt25BXHPVusQWQh7Wdgpthap+9dtQaVhL8EWdstNDgah2Uyp+8qKtWRG7
btPGXnC0wY6R0sgGu3qOuq6bQKP4dS3EvjuNpUTTdf8jH8GQjUhfqh3mZEDu2f+I
zW1v5l4u67CqZXjuEc2wUT8p+eS4losrlMM+le3G/rkrFl4ZvjmuZ0mOX0dD64H8
oWFFevT6a1GMCWTTosgmw9f879r4/iIKNJgcqj8eCduDa+XaUeW6UMgtej2/GvkS
s+RMcuMHSVLT9gqlh7UX2EuPOgTl6AlJHXuv24KXoQozS4SI2EoYEc7jpBKRuCKZ
sSpYPTVVikSxLPXEeX4DswkobtErRnlUFaRz/mCtDiXUKuGiLN+UL5SO2ZIE9YV9
s1Kk88gR/x8uoIHCceOl8E2i4ceUJhZbSPEK95xO9/79omRW5v7XyEdB+iEGPAnF
to3FvIhgaMS7fEal8m1fpwapQ+dKh+tRyHrVikmRFTl3e7L8QCPC3/3x3aaxjRxF
vs/sXQFX6g3/bK0XqKPhHxXMz6CYPjUvfA6JSbnU/BdZg3av7WnKKPlqES04y32A
6NETTu2+KVokGzWBVUsmMAET21Il0pBXCDhvxbVXreEK2pE2nNNu/aR9FrPpFIbl
znA6L9+Xu3EohYHLZmOVDeYSTU7DaDDH8VMdZA9CZsjmUvYbpPe+byE3HhY5c+iE
d1bkhJyjpkvcq2JJxvC9jEcW8EUynwmgbwwHH6AhRyYOulm70sUiL41TEu9LVJN6
ExKoObEVfQOzYbwritw9z4WtFHZlilmDG5HNuuzFNir+ER/wZ/9HkuFlK1lzxdpD
LL9mkIvzOLuThFxL8qjmNbpSlm3sHehfejeW0INyA9mF8YrpnNpTUUTqyN2g5S84
Jlv8f9nLCP7N/QyhhF8mepxkkqXJ31XXQMZBiDyvZyAnlxmLvC0xJf+I9p7F8a3G
fSKFVLzIfYik4CH0XPj8WljKXH6ZOIsGIWZJjHQ2HpPO6qztjV75ehccuj+oljoi
TI0Eu9wP8gWwRtUqgy5NkaQmyDzzXx9gpVrCxoM4NBHbjpDLbmQvXEQ8nZbYXZv/
3ew5JgpsR5EfTk+Atwq602yn5mWKJSizzE6bibMTVDXAFTJkBh0QAqJLU0cboFJV
BJ/jgVuWlBA7lV8s+nFXuJHe+JFmS0Nwy7sWfKX0OsYolpe7YF9XXSMLQ7mPA+kV
SPAbtnljK2jwO7Bex3ErRl5oIZT4AVTXUop4Yq7DAlvyd9Khdf+qE6rjOgMYjBWl
BSP+uMpM3JZWrYgtYbDrAcM6dxbcU/LAVxVYLCi0/Q5iJ2qBHZMr2tP5bflIJprV
yRht7Rh3yecd10VpnW+LuT0QglwYG9MGkesyEpwI/feL7h35/jhwebL+S0o0F3zo
jadTV8/1m3ORx4aInA8PSiABQh2ut6HrTpPp54F7OeUFtpMuibs1Hx3Vkf37a0CS
tO3faAnQV5TWfzGsH6iyh/4xdxzN0CSl2zyEu4zHN1mpQjD6LWDZqL/w3S5XsmHQ
1918lDyH4rGkqaQfkAY9UczvC174cdvbraknO+2eWFC5ByX0EdfQv2Y3f9xagJZz
1srn8HAGEs1AR+3Bo5JZP1Tl1gH4Vi424UOjHg1QnDBaeWYH0GrTt5SF/p5mU3T3
NI7LIm4+fiiLpjH1nuAAKuPvG3+MaSH/nDjKlxUTQdo43v8h5o3O1EDey6orFI47
O+rISCcLTasALmWs0QEDYEfgAUvivGOgCJQYmns2jbrQnpW5WHsq4JT9l6RtQYyJ
/wmRKIfu2Mh/iRJjJjeSs2ycBMh+9le2h9v/fF8TVCVr8OQ/NE7JzpzlImKQSaPf
bIQSNhiAv7kwU/EosdnKqcoWNLSSRYbLH03krimzok1WpfKhSSRb6dc3Ad0WIKlU
0vmtFBgwH+QpDICL0VnthtZcepXlJI/Y95H/9LsimfVOe9QOYWuduI1FCCsuiKiE
u+Y+A85+2v2Nq3ewaXdPlaaErlMvCN80lpYJHwef8Kpo2fjSmmW1LoD1Ckk8hTbw
+GDUZUgsCaS+CHt6yDtllkj5OVkWO0jt9IdvIkomWZbb1fYMXxTZT5JiKKOpr+7S
7M4VWOzZofOvcLAqDADiEE9ko8HYgVKjc7yUc1naHg1qWcVsEv4hRI43uv9CAd69
RPpWcU9lFCH9qWF8cvPCnIVTLpG8qMwyFGYSRvu7dEVAt05iJjX+YRmZ9HHU65dk
KLDoFUbYuCfNShOrbRbK80ZDSwI4/SUI96SNcKqgl5c56q7GliHaOZpQH6V43+Vg
A1Ak0dWNfSfznAKaAAOhjs7I/3hJOszDYgQ/QAYfZwQjQgLzzvCbjvvKGUw85Ei9
as4P7SO8QsEhkRrdvq6laKRsAfERSSAcNo7W68g9o0IgK85VKqs2qPKJSmE2zsRC
wdp1B4bnQzZRQDcTWmyN8VldDu/equuH2Jb3ks2RuPc50rTupLOjtZkqaAczra8W
2yB4OyycHV1pyPwppv0Bv2ioeUMTeRjQyQqfnLiOh2VooKZuQ79gUcVSVIjaiHZ/
VG2hlWhaiagLSWYnERDfPmPBBACcmFNXP5pqdsH9oPIEjgYlxpb6qT9KEPc6J9xt
KHkT/08OMoGDqMXTvMXo77gugyhYBnP2tuqZYsWYMEsLiKBk6L2IVMsUJYVxiZoK
FCkuMrqbsOLj1rg1Beao/cUJd24Joxygcz+bifjcY3qX7XTQjFE8u+nQ8IxYcHfm
dHIK+9HksjcP1LRy9lRwdlXQejanCukGcHgMV6+X1Q5pkABVhe1Bj8bpwuIA9Icc
jsZc7LEJdyfPmKRYuPKKXVKLwiMHDBTJyPbgeo6dgoAE4cGntpWNseI45NJYCja/
mzfExH1u1JOLm21DGYpu+oGaKY/wwGOVKAf0yVLHE2dR13kwD/mKL2gt8pdFOpOk
nR38LdPNQLz0zui80XsKEmxploFqL3HqlJdh+o3llw57sVg5g3HObXDEpsui2B1D
mFikd2Qb9L8WqNwnuDG4XP59ns0Cum7ZoaAOsPaVZOe1J1UDhxdNvsZ/FU43BzWC
svbad5wkUbNZvfDAKybd4MR4eoS40vQ97XYLRAksxPizuZM3DHtMZ+WqXMro/iZG
5Ve98y0kf7NN8Woq7B4VRxpG3r4YPbjYORCigs28HYZET3km7jHlFuqH6OXqa548
lSDid1oZKlM5SSVubJB1GvaNZWqyFbxp4BM+iaGfWuoq2FfYcX4BRIaNYSdYh97l
jKSyEtdr/vcxLD+nN1VUeyuC2+LFyqH3e9B1RZxOrrTogrYApDL3KIXk60KfpHpx
JZ3F8O/WML4Mu1NrKYAJsRciWUGPVQLyYjnMRz+KaA4gCMVDsVYWHcLm0IuyDuYs
2xp6Sj8mhQcIYY5sjdGPeiwK966cheImX9nfFrE82COn3NXDoBfekqpD2u2xLBDY
znnN1v5sU8D4wd5rLD9pR1/Ax55wFSg06RWk1TaEUsC0aRSy+h5Jev020ViY0eYw
Ti3SF8GwBvZZqTvsH2dQpLjkm3sgCYTFFCEG3qfCtUgENOXkvAyIHk+4LX9y98nU
6AOG1uwymPLWTKNtsK2sZGS0GsDoNwBAN7f/dCd2mlPZz9R6GbkzJzMLKhOuKpxu
u9uRd6EdfsehPGmX0DmfMhQjOVlmRfHbWgde6O8FrqkNoabWuJ5do3LoFNGowxST
55NzJJDzrC3ZXxhBG9ZOugi6OukfY/PH/8ihYw2rOSd2V0EI3y8LnQZ3euBKpFNO
oqdTGrAD9h+D8buFNnDKCngP6F2fiBovg4zdEUohdAZepYksfCzzW0CmTzoz3Fpy
eqBHyCxVRtAK2E+2L+dCjeycAWZv+qebSSW87cI89SadtWXLjXzsxXxX+t3PSrJ5
xpiBzEqe0/LdXlX2nOa01dhSlOMrVxlMilDeMdbuOsLRmOzivIYGFXS7Na3I+xKj
mCGJcrNp30nxF37wSIu2pzC4wByxR5NZ7xTVPdBw4sUuoUTaVE6/s+uAjQCoYNZE
X7YrrRrU9wY/hxzmIxi2r8CsluXnJnd8/asA2JGJYLizK/iYMG917u0PWbnwEd0X
nkxdnnvU1sck7uiQSnuac9S6GsjolF3x5JzS/aCh8atcXMN59b0DJ28ynxF33hm3
cc48maHdCI1AOkioLTb5u/0QE0qQRFRypwP3EVUzWjq7eTy65JyWxvOSnYDk8oBw
VzmmTaxKW0fiv5KPLV0CT6S322krDbXdnt4gO1cMGiHsPhKyIMGEVYfR23cZXKzr
1SlzbcNnJvb5G7sr0bmXIO+NhYRNpFNu9Z8RYGYBa0LSjac2IIGEo87xv2AKJpf9
vX4jyRckNwxVfb2Mg4pLaTcqsdOeo108AeWEoAlD84XQFBtZqmvLUd/cHS+/+oeT
vgdtmgSrxj9wkA2bHJ73jtUnAOpPEXwyD2739R7oYj4eBgO9TCiZoyiAKKPu6mjG
GfDYZ+a9s8dmXXpwo/Tm+4MSDL3T6H7qmKe7TDEpt+s60wS7UAIX4JSJBCQP6JWr
/N3UplVfon4kkMXe27qhEJHMAYsSXw2HQ/bz0D3WeUWz+RpaELNstCpJ+kYfNhsS
UHR5gr27leLORUJcSoPSZ0P4Ut5Yn2VXGoO3OhxIZS212efTPsw1bd3jmOJOFnPH
DuNio7fw/FJKV4jQ+z5bEClUXA3B2Rfr/zhQKF9bP/GujeFzv0bx4Kl0/Mrw53jo
CenSK9qYAn/oTZJZS9xca3QfExl7tgJwO4ePOawI47WRNr83TXbnT8VsXxuNwesU
rt73K5LrdFXApyLFHyXoyY2lgUZuoVDL8kRbub5P851Yvm+UcEhSbM62n/83gtnc
xmrIlTJoXvanJlcNpbSRzGk9wM6+7817LdQrTl7XqB2nTJ0wrD6G9ql7qnSZb8dc
SELFBwXeDALQZhQDJ80q1n+ecCfVmxsinuM4IHVef1v24PYgAF/z1lbXHLu1HHDn
/M+7FcpGXhFmyc4lSazjCixUX1NQnINZPZAyNHnOj+Z9EnBAoOziHYZuQThUz0kn
STU5puDPNxmWN0b3PySbqcQ0oFv6DeorhIn0xw2VHqzm7TNHtF4XXvUt3Qx47SwY
TIb9DeNkHOMuEzZnOMZvIVf6xnV9gxUOW1XBk4V+7lyndFBxdnBI6e4ElOI4Hvra
YcwaNO7xzL004gOO572jd+uwxSCgLN7EDtdCJfokMGX/VGB66BrE13ZatHxxwIFe
287FOOkx7kTkov2nCqk2+kZ0PWsbbMcVAOM6Tb2HBBGJJWhML0fAIlrRNj+VqftB
hjXy9rPr5/KInt3Rgnhn8PUrqXR1KOOrg1k0s7RprFEbI6NzRMjVWQUag+VOqths
Nbhzjt2TfckUi4ohF1Oj5J0yahHqtXYstMhUuIedlTev3dJ/9PkRTPwOng0NY5WY
9bHQuzA3Wc5uVi13VCp7jzLvGrUXebRHG5nVq1JqFze4B34mmVszibOBQvCgfrxl
IqJoi0IfsqLIEO8SMSX4cU2s0n90crZrPFm5jhfYlszTh8SfXniiIsJ+LsVZM/AG
1qQBN7erGf17i6i9JsukXAcA/M1iYbHvOPdeuOTLgEHC2zUwNP/VItTGFOuo5vcx
loSdB5OHQ3aNw2OtrrHSdiqE/UMudLnRUzal7ids78+/8OYtKhT2N0kPu5cOX4yU
rbgaImOra0XDnhaBOAfeoatUrgyt1Jsv3lQbd0xHjkggGyH0DGQLcxubOiR3tSBw
DNxpsSuB2Ig4j3tCHWvKBRwU5JYhvpfz9epl0Ss2jldbjYF3My4L0MZXR1PNRmQ+
n77kt9w47SU4VbUMxIEmprOKdQJY2uiXSmi2q6dGt+dssdLoyUA2wrw3eoiHOb7/
o6NzHvWORz7BUJA92QM/Vc71/Pu6ZfXOR4zXiAEW5H+WXTfya9tT4xsWkgr5BBSs
fmk4q7gHw/dhYgkclUvyaU/xZFbzr2ArH9XhARdc5O/ZcnalScmU7HLc1wsRLiWu
iRkQ30kB755kADwgvW63WYTHlt+UXIfovH70eQvRwqZW1lr0sFhjSbjhL/F5dSJU
7iCHDnDYDoEgqahP3Zd4bD7grrCC6bycO5UUGcjVjXHI9hgV0Z7Pn0dpm411sbIs
GC8NbWMbq+Jqcp6DTWMyijypoxs4OIWEDeg6yOvSgjbZO5m9uCRIQvCxbwvlCDu9
2Xpr6kAHicNAV98yclPG+iA29WnZLk65/Afv9o4daXHMXCA7L9SPblmv7IUl87s6
su0f+VtQfOKIJQGzKcRYP7HU6Pgon8LS1xbjsVh+292a//Y9xvkUwjl4r6bnVOiE
qetuLuD0SFs20eXFmk03RjiXf494eRjcygJP1Ss6AlERA3SWJN+sHT1CYtqClt4J
5KNcP5BOE4Cj9sqp0n1stZgvkgGBHys6MSmSAAtL9o8jcQkJb7Y5sWpIzHI7UUqV
VwNuyT8SJwQ+xrDoxoZeInbkWk6IF7ClYaw9xW6DGBW5m1FQfNZp9XF20v2pwh5m
pFJSXTkVOq+XrnUNToHGfDjqx1bGdB3zzvFv3Rn4yozSQQGhK0VC6irP2tImc6zV
ZuDv0JKOuEuMu7FzQcXDqtRANERPhPZOJ16jhiGjDzzP/UyLJ35Sz87Ka65282P5
ZfgJXu3yMJBrkxcLDs1hEJPRuK6N1vf2wvSeugojbayo356P7m6Nl5JaBkeLnkaL
61CxU+4UwM4VwctDbQcqEVknWAadL4WOnGLwYB8UAO1xyfrDMLilxrqxyHP90x5h
Wl+bK2Jgd+r2MFifoZWvzYJYN3VN8mMzjf+1OtaPUrmf4W4FyqJNXZGDBaDJyrjD
mj4/Z/l1I7jBjsaiV9qLO4MgwVxwyf7q2G3KUb+Bg9M80dbPICYLqHC+ACA0DtzG
HemPL4IzsBx/auwIFtwOTRhJl+v2NQpQtYiN3vAnW4D2sBhosOcmuzAWM5oVPeTz
kYLO3lZbcQPEMHXtKac3T1c1tcIEKYPk/jULQMehVBurd0i0gXHDy8Hel4oWUmWy
2aps9d1zVPRmhouPOi658nD9SbNFd+y/9H5GiR8JVokPskyo005RB7RHtGtPn3ii
0Mw/sMm+1Kmw9y70/IbYpVgAFrhJqCXcjp6f2an9PkKl6gnMU6O64maJbEenpJQj
CFSgda00cwDxdKlwwnAmaOtGwaWyicSc7sSlGzwxFvOGwcBFPt32gGy5cDLxZbl0
Z/1FdW8MM7p/8CSLb84thuIPbdWcPHA7ki3iu3gm5naNFkbqywKyupBauDzK/9Is
+1UGY4fZEsyNvv9MZ4uM6pyY/ni0eoCdc9leU/T2yYCQCqxNiIMW1GxfCbL8bIwe
gUktMmoDJg+aNrLHAvC2bm26wVJgtkVeoQcFLojyiKE+05ddeepGFTFiQTBdTDQO
XeVrc4jS4RbwBl8mPzDnOglTYv6qWjcl6liY6PlNRx4aXLo4MHAbJhwa3q/noW1R
it7E5rmWPhOE3xxhuF1EpwI5r+LOq+XfjJfHUl6Kzya0SQqJrhbbukSyFYMnKIdK
2fiQ51cYb7ouQC2d5VufUWFtGZS43lGKDAy4py1wE5Ixsqpx8GXmYU/BcViTzCpY
UxIcEXpEj4hFc4oMtJc3pDY/sDrCnYpKKousdpUDjFMR8wH8jxm7DGEJIAVte8Ex
jyoG8t7P8fM6kZMrk81y8RLwp/gPHTV0G3QIkJUuox5TVq13zYpO3Ern6nMErAqg
mCF373SUVBK+sPnLyE+nLWPUh15ym8RQhBxsrk3jk+xBdQMyPcMczauxFVfEp6Tm
r+pq6mw0wkt//n+A48OkGbYaaskxzVW+plbnWAcPX0f5hs/Xu2b0vcdZxmu5U/sd
JvDizlXU3KZjSRSOSOBr5GIXru/srukNvJB9LDpqZWDu1Em+0Tgvz6K6HH5KXUlA
51ThOjvPLvcQqhh9dz/IpsdCHx1htXKhQez6KkKPgIAj1doVxMvfhtx2t7AVtWBL
LaaBPACuMoJH1UrkBw4GRZUFXWbNr4Rc2BRIzzv25tWOUSrnT70UcUdfkMjJw3rp
g919pf/bzUdO26DJ0jxpKuQsXrlMHENhF3so/JmPNFu/mq/MGYdfLRN9nrZGz0LL
78K6Lth5tUBkszLhG5EELCouFe+sUwd7hnSWqFAIjbSeiGk25I/VLbQ3AXCoYwlO
MsaEpf04y6qfkhuDIe66R7ZPxtP1l5lZCfBE2RR7Sp4TTdcj2Iu48NnnvmJPjt9P
jQhqYWBMO5HQ2KqQ9NtIsup+FRrvSya+VFj65AkIiDHPxUOw1px2t09bXpHsQwe+
TfYMm56D1DrPsXz6boc5nrRbAgH9Z/+HuCVndnm8v59BslYoA4x+k9BQJOta5JVG
E2K4SXooYoshedJW8WOTGhX1ZdZ+cjHMdmOrmlztSF6wOZZ8NB6RqsirZ9XY+N/8
QPzHijuJj4leLwqjCqiYpgK28kZ90AliN0I/N8P+kFg+KBjFEGl+MZ7yGbF+S9dC
+iHBeLjjG0n7Us1wANfHvFti/PvTZ2+ojx8k5c7qT9Ar1J9x9nNkG2mtvD3ZJBT7
7Va+07JhkYoRNqAGMlsqRmoqPW7wGpMdaza2PRJORw2xNbBWpBbPC3r8SkWTIiSe
HVMfjWoZNgxFcvQwkwPaLF+sXO4cthVkRVvVIq9Xyc+mozTQz5i4aZscrxww8RXK
qvN93JKggVY5r3Tl80yGDFmiayegKX8KnqVDBYw4I3j8ftyesmnUCkRwP/8KZWGe
gnnwAVKVBGwjdalGgIqLqEM5Zq20y5Vk/Tdkztbwnc1X7qyVhfGPPUHSur/ubDrc
RW+/WGk+a89neMO58xuWNl8p+w9DCIiSkzG6SfU2lgCOd/A0Qg61j+/LpiXui+tu
5trIMi4nOJYiffcGLk3RXML7UAr6ieNYon3FKoCxMUtrUnbph8EXfLje0xomqOHe
gABv92Jmbs+z0otjsei6UYjHDui6rMeAXwrOQXC5i6n+69mQtQzd7gaEOdIa04N4
IS+IO4qEkEfo9NjG25vrPjfs5YlLXPN64Vzn+FpsZOAN95qjcN/zGgvXDLgu5mDw
ZZ6ruTg/Zki3XpeLocpSXU0/2kpSOXINlHt+oo1g66BFXrAVGJi3+YpI485YRoFY
UTIyqip0EJ9Qis1FfeeyJsQLuLBD3fXwxoKtS7xt+o5x1g9STsSRq2qPIDXmOc4L
+vlJKmN1D8SvUCQGx1/Yxa3+sZkSrL8sjSFBZ8M9kRfFNuXgAs5IpMGI5Dvzu6x5
a5jg9VKb7rTKMJGz5/fBznDOcsE+n8xgXSUceg8JQ3wUEqNoc7RHz6/SZv+Ym4yD
wbkzVAugCDZEwdZiAgXumQ+uBVYNxtkkqBlyWOKA1XOF4uPQ/j0Za9AAnijOzo3U
8NF8vD45w5cMXW8/Eog196UyWBqansAYFJ1LQtu70wbmub3D5Drna71sc3mHk7Tw
hNuNldxHkYvFPrf+IVRgBvhb44zQy5NWPiv8KFkfPgsAuEFNRc9JEfSIn0r/DMCw
AcYpIWOd192xfRqrVK3ia/EJbS4WjbStTEdDF6JHyC158bvBTmaLRRp7D+SimyG+
l9YS1pHN7eCyDz5309znt+lWgC9TyZIEF9I1G07x6M87swGqe2F4iTY3PpICcokR
iQ1ddpVCI5kiApXoxKKLCMXcCLJvXH/YBK429FuYG1rYdGyKTUHbje4NOMZLo7TA
jwZyufKKrVr/P1+H2nVuUKQkiH7ynnDR5CxS1Ou0WYdMNH3CLN1XTfMcpPqAcJuk
WgUntSTchzXFYfXaDdtG+HAOPd/i1w7yf/3atdZAdxfKGvQQYKLHTnp2zvXjrdWz
rC29Acor11s+or2mpH8kXOQAaJHKv1LsycKiz/DokSGqgMc+DcCNc2x3ndUJG/wL
wJKgDv7Wuqd8Dzxf/c+OGO5fjaL7x6QC6YbcNtgd2YgNRWE5hPm32fksMo+lVhib
cesomEKsXHhW+TNjgMVr4KNdtgh0d0zUwMyswCCezWo5hdskMI8B7vuPaTPI3WCl
vhmtgJmR2D//NImQxr7bZdGjWAwMpRPslbAkIyGALqVZxIBhU3zVXWZTRWZ3Mm2S
YwkouL0+D7txqery/9UTwVZVM+ugF40Sejxp5W12cfm+K/8BgGs0OxjqrQzq9lAj
F7LHOQrbKMcYGH+18jMblSqk2R5nTNrJOUv5RNunUfrAl4j1DkTvvNVK9GQZXsqP
FB9M/ETwcrTbWB+CUg3uFzLxgFS6CVIjVVXPZe6oLCT7UO4ZLZDrfZt89e0nDoqO
2g6oJGC6u1QtQyD8L/QvXFSRUpdCC/W1m7CUWzN30YO8Thfjeo13tbY+AYgp9laj
4yulSr539krj1dpwh3pvyUQAAIrJFvV7gH7ZCa6ZATV8sBIoH4YF17fqK/X9lbfx
KzrOx5vAGvwlaYECx1J+0M34KMOHn5Cxv4GdB2yL4ioJw8GDISek3tDBB6PdF20N
wbBTfDdxvNNyGjznEq8tQvjaJUgt9GvLj+FWt/+VYpYdTi+jnpDulIqS85XujVZX
tKDNXTSiYl1IsEwYol0MwOEJgsM0GTv0roTJ0hx3DZ4oxJ5IgdgJAu0lnSjg71jL
7TvsuX46wEVxlz6kM0pSeRZn2gcptTQqsT7ZUen8wPPzzNMhSyYqZqnTXyEGyShD
e4ZJ9B0X+Nj9mmU725+QsoJpzewGbAFnVRv4Z/pc3/SrTN4YHLbWjUbOzxNfBnmB
onmQ3IjSYfADtmhShxt7r77+yHtfqKupE2p3YrD/Dp3lv3lInDkJFQ0LowWP2t94
us1E3DPhltwTPIKeEz6BJtLtNLsXdy9XKL6b1Rr5e2042cQSAMa0j7zug6r/aWD4
40O2deDZiTdliHnSvOh3bs1WRl9hl6NJhiYkN/c5/n09VDoD9+yjx8FP7eliAQzl
wxfajh1qdptqkxGyy2A55qRPUXuuUDnXOs07ftiolO6z96WhoQWhL4pXjX7+4yc/
7C5gW8He1FxtJJ25HUF46ZSAukGejw9U/dKARp5RX+dTjEPfHZUDPECG6xPMm6fR
6gzWfzqXuyRYsTHwLU0IVHQD8ULPTyAPy+Jxo5yxRXNXDLIBvWM2pDAiiIrsUJp9
KeSE4y378ClQPV3OjMbnFNWvFTmMPfINEbsyypYhjEOeJ50DXvKkiECbvoU/7HeD
sxtVlRaBjVix2tgDniTeQQfJetIkPaI0y4JMjy1GHTYtwsMGv4Dx9o/k/KmHQ9Rt
t7r7GxisxUIZDEhiYHXV7b0BfoZV9Ct9BqeEUZiUVrs8bvho92BqZELgQBumpC/i
ngA4OE299Rq9sPKeweQpRAMdQiQ6rfljXpMMfxfat0pByTSaWlnE2zy4vWMR7+oX
fdEAbLAx5ei1OtJKfD98qM0o5YQJ/9yqEqCEoJR2qP164QUhXIeRqB2uL7BIgXxe
Lcbd7Tt7k1o6IwSsFlbuFCYG+OQ1k1rpEvs9toI4aaCna3+FgCCevWLfh8NiA2tI
INEDyrgvKNNjxf1tVtvrDYU4ByDJEu2s1YxUpJO7PSeIts5R590Hz7Zcs6raODSv
wDflcLmB833uqea74opWfAzjKPB8nJqRnOtM71nmnmZah6JKngPD/EfVF7sZgZ+h
HfnB0Zo/2MW3z9FyVBUi4pMV9vJIdLEZL92u9zkgccIveKJNhbKGwc6d9g4Nhm5q
cyb5mVCjqSnWQgAz5pe05VdZIDW8ws/IJ3KD8Fo4AbAuOc3Zn7MXWvcsycLcOzs+
aXLCb4mXCmsaMTmaXtqzVPqWxwIOpCWnJMl5uuuyLw7wRbB4seu/6Umu4Lg8jUNd
z9k68YLGNinMGHWZJv4lC9GfunjKAD2pikmRZEQbkfFyMjFuAwIQ6VLN4N3R8fWz
1BGNhH/sZOxR6bmbMJhfWwJCd3S8fiv4XJLupHuTuMhaOPscyC4FTLLlmN5mflhd
dLO7c+9GrzUBtANnhiPWZ04WUSJpXuhQgn3FYhLev/YNdBGswmMUh+FZt7vcyvLy
A0LA/JPnEM2XpIbCLkPic7lP1+WfIJNEVyW6JD77PhcpoNQ+0epF8hItJu7CP1AS
/jqdgVjIEYjyTgPODD538X1GkTuvAe0ZWFvDjctN9n2dOCioOF+GUNj5k/O4I+Ou
LLGNWMdSGHGSnce362uY5K2Yuc09cdpM/q88xEl51KvxAC5Dun0hqRcNDAgVOdAU
7sLrixgA8ZhvSLuyoTFSkS/B+rHpH3X5+BKAHKqYROx7Tiv2NiqZXORZcRnZWl11
w1x1HbFCNs05f1kR+ORO4QlDTIOrurysZLDCRsNiRKOmh2xoqsPSi5tVLepZtyYD
lv181hpTEPINHrjvc8bXKaUNaVhp5DdWT7mUlguXMLp2Mn1qGYwWbmMLQx8YVNlc
xCUuul6n3NY1qHvgJE4naVxMAWLoilGi65VSA/deK1uVghVENPQLO/G2UtyJymFm
i+d+99dqJew8hhHs3uk47ddiV1OOHcwWB6ggwp8eA8A4GqAby9hwbxdx9Bt0zwaJ
f/Q173t0H2gFxnaFwp3tZk+OBskZrz1GafLQad5Z3Qms7t2xtqDwC1Rl7hwXRuPg
qBEzcuhXHtb0VU1YtMZI7oB4/J+HWoD7FJeXiAyrOxiDz8muFtrWIyNqcF+wsd5Y
mdgnHQ8HuSnWUcdbCeyr9LumUw9YoHtwLGPW0iww88hla8Q/wF4YUYtN8iWcsnJZ
2p1nUtcSyQLvJPY/JYRe5lEkLCepxoz9Tde/pP7HRU37oHN0h9H/YeUSAgV4dOwo
P/pSixR75ffKe5Qp7whgoaoMzqvQax90OhkPBGGIkFOKmjd1KYBAViAE7ek52Rwe
GYu8lgETtvonQcrNlt8eNekjrmnhUyWanEoW3m0Uw2PAGFN/9P9J48q9K9rgz/6L
wG562k60wflXCc5sR4+KiL6+u3iIIP4m6wQ/iCzMZ62rGF+ErrPDypoSHabWFxDz
jqq1+pDIBpVfS1T/XGccRFNwjEF23O90QpWSAvr8Tyc/0LcYpHL/eLhaQyYg3ExE
tkZGptrwfzZlbnVo1BXluXiIlfAq/dgBsmCWM5EntT8HYhIeuENIVBaQRYyupHS+
fsEnr/OS7j/JLxT0DNLm2l4ARC+/77oBsbyC6Yc4IcXOJa7WfQvr2DUTcIpTIYLI
IH+8UBsJddaRlMYNomgYiqykF286jm3ZNGA5U8Gebb4TLlZwPPtTzdKMoGX8PQwr
jeoR+fSX/cLcimFN+Q6PcSCOX3eq8xI+QMxHWstMRETcGqGnPdm8OdWRBNh/uRxa
zDv8Gor55GbwbrjRN60uU3T+SiZAsxzyksHLm3nv44TV2S6CYQjyWOt1diCQJSs/
J3C/A45Z8OEVV4ErLf661dXHcTEYWCnNfT2OpIPRQ06/aKTA77U8hGd5I5HQmQH/
w71jipnK5JYDse7hMtCh3Nxo3URZd3W2jd9GXL5xlFsojBuAHGdWuKeHocf/lPFC
OL8C0Y/BkMQ2anHWoFvuS6NGJCBFG8y70K1CQQxoXb8Wie0wTBvUcwQSFhu1CJvI
1TAurFjCL9mCYNvhqB9OsMc+FEfbvwm3phTYpBjc5tSI5qywt+ReMtUcfI7iuZ0w
4A2X8nmQwfjPnGE10GxB8ZPG/fAeA9n5PHKyqbGKZLNo1/ZzQNhLJArJ9vz6lM8D
NHuFTdup2F5kkmQpb4SntE95WiCb2IMxtY3Iteen4Kq/UnoHe/wq6e7oYFo6woHA
ne6NF6KryodHafn55UN/FW9tR/hhU1geACo5COn1Xmp6EiBBPC5c8R7IVt1Mgfel
Td73G2SuBNjOshmME7dfe2J+oI5aMzw2yvgpZ15xGgq9oZF21ClDwyXmkFf9egtZ
GPbCubAQCLuvahMxb9/xPAEqLovmiQ/M5E8NkB0oq+oW6NhF8Zm/YP120Y2EIZKN
ZkHUqoxQBdMGv7iBzPYj9MnCh+IqGeRUEa17vuLO5GhKCICVmZXfdvB+SFrq4tpe
zadhBGS8MxPfn28h57KsIldn1EBeEIpiZ6wakntZXF9U+rKXRD415AdAeV05nUbK
DH2byd9G91qTBspu+7zwmFXksrbIkDV+KNtGEn0QpOaYLNHyYJ247oNHXdXftgmT
a4nojuLfNljWYdRzmykDFZFnqNpv2ld8gPwEkPzGRFD+LhONdvzSsTtOeYdg3K8S
tlq3YsRrZlNK8dfobrFdfRGORWfmGcmpJvcSnkAyinB+duatokp+NjbTMByMQWmI
AL0bsIkznYChMHrWPSwdEXnNj3uauyMAWzeVMjfECTHneT9LLRXbp+XvLq1NvgLG
Bx7P8OY0Uois9YIK1RQHN2jDthgkED65Tnwt2lhHkZAKQZNjNwfCdegqIikxWkb4
jhzFXwSkJoEMnqTYx8BSDnLflGoY5UFObIyou+pEOAfNozi9tkyuo3GmvNPXplPu
qwJ+Ny4CH3thhJRVbI3lxb6scECV+PfBtvTQvVFqlgqAhX8Zuywx+L0ApDhyeG1R
IBvJ/KoIjB4T4K5+R5A1rlQancswAI6y/1AbU4NdzT7vG6tbceuFNitfLeAvgu8N
QFGbfPZeyvazBGff7hG91DkyhnbB4pdCLtzJbPcIyUXrFy/ye3N0+pjXeItSa6wz
4rDQbYFhKPhPvKQ5s3ulsnvgQXmPITxqWhdSPMdCbwdPPso/7eNHrVF+vVYBF6vD
p6FOysWiLjeNj511FopSTT70QiYuoZMYtCbcJN8MR0hKc98PbmNQM8epIN2+MiBe
xhSF3ymlWJIPRLxDI5jUqwl17NXGeWKLE5uhbLXvl+dAk1IRdXPzc1Bt8tnzsUo7
+eE/JSPY2mFLvecoaamLPRBKDVl58PNw7OyzMyW9wUvAKXEeXWFYuJUW5ev+Xv9f
2pBylY/Kn6wDuti1dYFjbAR9mamnlDFeidzIje6V5rYeIS+CY5u6onMBsRA7QTwO
ko5XELZ6TMLAWQwF7d3z4MaL350Rh54eozkZGp4gmyMza8gopoXWnX6ECeuyTMtN
EUMY+WO6nzSyPxFxjqQsfEtkmMVsrUzBEPeIqnDUaqNGjNa6IgcTpGPEKfKJtv3v
q3DM3C2btM1Q8bBN0rNOnZv+Sd6JLGLbb/WAN9vSGNww7mGUupsj8JhUBpE8Yrf0
ZfDiQfvGRr44odqMxW13o3mJesypThd4kZjjsc+DZu16/hXUGa9LaGEmpd25RfPg
VfsMDvwq9XusErSjYF7nffCmz7XP423me+GgdXmadRArUarqlH8l+xKflOnx3Iih
OGbBp+rg2J6744zVvIn48q3srCvNlUm8gw1wMZsyfZSLgCftaUTtDd4LF83RaUSB
eYGVhvdHm9+rpOvtIgd4CPzopYw0pNNtM0FYj6BGpvcqxgGj0R+0Cyh9hoIhnETC
Z9gAgQHH1EXcWbaZpbdmB076M8QyizMNDnlO8jWDoLlKzLcdaC/TybgGzoUCHSKw
m08PK8VmjobXVfZQ6pjApqR3KvO/gufzi2POw2gqleaFg5M4sbXV80kR4MdNmVbG
p2AqtUUseuK9zMedqmWEy9musf5fm5uukS2qLCHvsMwYOm2CYqjfGnVMfbU+ga8q
QluTy+X3aFK66B3gCb+6OgLHRqM5C39xjiEtIdmg3/1nEMF4gNVS7CTSmpDdYqfX
sxQ1OIa5FXLspFg4uMYyBDlUCtXq1Ny6dGyt3Xw8Uw9K98rGRlUTA17wGfzpeL+J
fHecKOwnG1DuzJG6kHZWVizuiZHtOn8lGJZ1G43E8NXXdlJCRu+GaRB2tm9Gx/e7
FigEaIvywA01tovbWiVjD8QPkC9iDxc3aplhYnxI8c3rnw/zpt6kK61jDRQIVRPE
cgyN4q3wd1AYNo2ESoxtheCwWTV3z5aZOrr2PGRHS38UYF1VEBoPGrrW1paRKfZH
NA2dO3Ti/Vt0eevh/H6zOjSkW1vbcKkHG0K4rnAOWuarxtc4CwGsb/2zrs0d4VKK
/JzYbhrV98zP7B+Kg3jQmmxeYpzmNmMIIcBHWeAA86aQFOa/DT4P2uRxIlvJi+iN
mpfkcEDhjiZy6fLPRrjYisR+INKo9C047dc1PMUQw5rMzEWThW5yM1R0qUwyxT0v
QhGiG2EMOzzVF72qUYysVWpHIFHJ6mfDL/H6l1Ynw/C5v5wrPYpDlGlHlXQZviGP
fBgEdrE6xvmlpMF5Cin56dsiah5rFTKTuH6zq2uRWNhseY2jUgvkrIdcxOwAAWdc
GJWWKY8gJ83A58LoKKhPvlv8omKY9b6BeaQEawfBDK8WFtOTbiUwHZJBaVFx5M8/
kXPsC63SxppbBO94YgRYVguj4HK9JDJ/HIVfPYi5vpco4ZdX4H+RyjTX4Ih0Y/3/
anStD2+MD7glo/W0EJ6pMzB9K6oQXrdueCeebGAdo5hjHsdO3AdzL+qK7xXO4FIi
e9/uCFbw8c3SdxWJIgoZ6XS2egPd3agL9FiakS2OsAi1IYDs/+30dGzflnKUzphS
wUS7sK5cvmHpcuvJT1wy+DYjh5/HQvCCwFgQdcYN3r/80CzuEbsWCgBQMwlzWB7k
wGvW6Mw42Lxa38hxk4TTxgfBgkoM0xvpwd2rmd9gG+jVBaQnTZf9lh7wvqois3Cg
tknlFqznQoEnQlObiC/RS5Ir/XFwYprYPytZqizlk3K+8I9avezbtX+n8NPxnsiq
wL/hLrOzn3k2BhEZbLZJg04FHAhkKLI1DTtW6iPo0fhvNxBGQkckheujRj3R+dcf
MVAquXL1MfK9pX23BadJ5eCMDrDNMTttaO1BS5R6MXk7fvP85ma4wv3eJe1wg/QO
iTrZ5lqB+RBLCHKaDBZG7yl6iwnD8SkzKzYtfwwj4Js171naJu6oa99N5ShwRBP0
xFOKYmPnCaotUew5L9pxm9sFAInMWE54ahjzCuKWAe0DQ6IIqUw7Tfedmg+4FhfZ
xXLTCwrlbFastiRpmC5zbztulWObBynBgSz87iz7H3SF0y7LHt6MFeOI4ToI3lnR
lld5xXSkZxAbDxLZ+umLm7QoQxqObCl+2WYHcJor5eFkCXC3n4C52JhgiYmfgvvB
AXR2I5Xsm+s84GUcFNhZnRkQNd8jsIUhakGOMU2NXPixssAKD5xoiQEf+vBEhPX+
o6JE0QGzgPzUNhHT6ocOFqc2eLWfu1Plfegu1fkN5RJ3O5O/3W4f+gKKHDZ8Dzt/
RZko//Zjq0jahEc1cPJTgknPaKqa0aDzKwF5sFTdTvE4kqKztAOOW/QPoqZeiEaf
kP3/oyrfpLBJmXGkgL7KiICT0wERUj+p2u2hiC81wZ1yMYFtNaLzC46VveOOMG8n
YMS7ZGsP6ZC3SIYpaTZPr/UQrXc50GmYYSLAhuwqCRgz05ZVV8Nbp561L4SLuzkM
Sc6zIKFjKawwE7uWFkyELPH1+5D1FOoti33nMwJtcNIxFLkbSEnHPbRxziEuuZTy
LMQuRQQfoImkFVZmpWeAZfZ7Y05BS/GaNWm1QgYikLeXKHimP7wjsAVqrmxhNwCc
Yh+7O5NeTIhW9mmtijiz+T5v/Lq7uM2ND+Y1j6ZBlmSAn51pXBpJmODpjtvPKxCl
+7Mcax3Thrn7eF53JtSp7ywmRKnxzZ0Bn49GDH7fqjHHagpaGIbFxGmuvLriHodc
XW7AJTfAJgqahPFG4ssTF67EwsE8Kmc6NZUgnZLtH0mi50N3lH1twS9GPdK0ALK/
hv26eu+Te88+j71fe20awbVXD0J6RHX1iHzg5lpITmRoF080e5e/HSpV1v4m9LSa
GuVo6exnDmKlyioTfeUK6ARIWtfAWk69TxYo+drv8ZG1b9g0C0ZFt4Qtktj5l1ku
VviOkLSdflM2dpjciYYDOR3Vgf/am0C3RZ4e3AdLAl6fZoQMJkS2dHyHo5ivigyl
VgpTWYJAKJWRPm2J85DFuNvshjBwnM40adrtaxmMYAEnlwjsEi9bZRrEHm8tV+8Z
5XvJW+HKbL3VBxceSVdcLY1t5NWIVB3wnILInp0VNKcI2UarZU517zlq4lRSc+kM
RKxNianyTSuaFvzHrqbTbFkRHOA0E6gcoiaP/b6LkFq7+mj+lJCLuMwXt/9xid65
+OS6ymxxXt/+nd97Ion2q63UcyTmELsyGFBJCDQu339Xz4rCd4Ai+dW4ZN5a2AS+
HquUsi0C4KhJDbVvyPkmkgH7hISbiBS7+m6Im4g3utYYI4vX/wnZpgmdE39ceoPn
Gm/uYPvuYGxPFxiYp9AmQMphZJn9oZdx1m4z9/6DsZygukOQbGgm++LDJYJY4WK1
Jm3Z3BejqsWIdoQadxiG2yQ2SWbTKv4SMU0mLRhSpAgqgoC3cgj6O/HRFw0uWEDj
njsYe7UNNPtFgWwPRlDMN0EGcOo/4rILqhN0daB/3W3UieJFXqTMP86t/SZLxLL4
6qrEsHw6ZEFhTZjtOJRNM7n1/J8XxEs+9HiQGsk1ojhtqTGyJgvas3et/xV/22kS
txW2BUUF0lcHB10252cyV+bbBi4mmvbXbYuzUSoq9xqZeFh0olGHBWX1dcK2f7V5
vl2TjZIza5QIQB6iEzECib2dORLqylHXPvEthTme530l6GThaAbroPboaFM9jfoj
8ZInS28qJNNQSk1jN+d966Ew7SH/K02IGcel5Nqu5MhfWuc+ekrfMURdYEKhXfiI
OPsmPmhYcmqGCbsUKzrb8CetfW3MJon8smDx0n/vsbQWG418jSuzx3Yr901Ha+7O
2PwGkGlB8QIccFZ7/LbrdS77g4hoESSpnyE/Z3LKmQdcvbIC8trVb1FY0/bsyYDm
8x+12POt/QNFWP0kisOl6ptf2kpX4QOlwFy8V/dk0rwrnzM2PCD7A0BwUZTH7VZR
ZnicrS6RECRH/DahNRGYPJh+1h5dA2CFQR70dss1+WZTPzn2rr/gYtWMGAF2XduZ
U35nVN24GGx/Zd30CZH1sfwNm1A/Pgb2rQ2WPEFLAlZIcUg9EC1T0uaOhSCnG1Xn
oazYMgLpccxBP+zfeCg5gE5e100glj/D5n26CanG3befXe0Lu3LzFxo3EIwh4Cd9
bFu9vpY+nX3cGmSm+jScIrMInfTYSmfv3yrdV2tiKzMbgu4/P3fZp/tZbDgnVYjI
hYKIyuWqUq1lwTOjqbCQNLqhUuQUdOVeLEoEgsWkaLv5u4Pc/aA6QTj4VErz6Vag
88c30HoCjw2JsfbGA/RQ9HFgVXNjGgUE7YZDhe0tB+tKQgBXvQhMtvd469z05OSV
NGT0466ll63hL1/SE4gIfV8MczHVfDmwDY4pv0fkfMjybcYuI6L1wNYnCycBQEPQ
3IbN6C8tpUAhX9qNff0JVRlstMZIEJJPWTGDsWP7Z7EWAYzaKPtGkHfiKwz3rtnN
TGoGpNipmyBYik94W3xhjH3A8keMwUuQYk42ix/CZWHM/ovjGEotyYqcL4aUsZW3
OGUTzp+bDb6TU+yUvgwDdokKzewJbRPO7weXkACB/NsKI3wTNA7nxx2v2x+7nG5T
rSaKUsDTaBRW9JMeTW2eWQmsyb2EHlGLdo5gBA4ZgWSgwWXsbiEErjdjn+827bZ7
ClwTpHlTMOkCU1V4R7+FPc7pmBcXy9zQukrWY8paFkuBJaxyTj5ZQNrCIp+Jql+j
WMxg81vJg81y3T7PZc9gSN/ocK+VlmOllbcwcdpnM7sf7Rob+W+/UibMXi7VFncQ
8bOWRwrxJitAiEsQ0kHPKlGNTFdiSP/lQ0EJE6F9i+y7Wsu8GzaCQ4uBj5WNpvwM
06w1idjVCFtMpLVKuHA+XCBLuzXV0N4+syMRfHp6Tbt5B7ps2yUxAvOvOZlRfD17
KPxyvBy+niFp8TJ4dHC5JrTsVv9CurqcWXtrdtyqHYZ3ghpq5n8zFQd3m4DbRuIt
OUz08N+Mu/ednHqBmHkHXu7qlmnlyweYvWhIBhmBXdemUop1eRKHQCzR+VUBsXr+
mJO13TArt3foBO5qX5ZDUYYifQin0r2rgbuLaGqDq10EMNPnAVxmykNd5ZSG9Uwm
swf0K2aff+/SiD2UlH3hLPA3XlLJSy9VOsQRV0KTgKFpv7O9Mtz5HeUjBx2Z1V5G
f6C0AOAlCZu11ctckDyxLjTcuUdmfPmByztUd5HjqS48UY+8ZHBfxGi6AigU37zV
LYW1e4gUqGe08d564VMc1LEuPGRnZeZbB8Tz5JGgoYkKrVjPCMKwJ9dBaqkjlQJC
XmLtJ/rcY5P3DWxEu1qIO3dybXzsVqQ6Auk9WHTRiZ7azIyMwdkNDBf7v8xHXLbn
ikWNHeJfrk/RMc+R7d5KZmFhCs/Z75bCyaEQH228jcR6eP6jSySZltREYp0xdjCR
hgNLHQH4+m7eGopty2NjkG1SNwvwBM9fLDUQTmYRWvP9QGBjjL5mNcgwaqfpMeX3
nLXkzR1RQLG+8sRyqCMMmg3sLmLRx8yAb3S1HHhBIppOdDRRh7LktolHH3qfGiEJ
dsfEsZBLS40XntwMALtcqanelCS8dzPG5EXE9BqoRf47OyqcXmiPAMVid6sJKOEg
ZwBnkoVy4wxouweXioFzlF3k01VPj5ungl05SMGTG0gz0+UkSRwbE04P6um0MiKN
RW2a1HU5U4lBDDT9ZzF9UuP20bB8LdiuLP9LlT1wfbIuoeeX/cvwFvZr0M8GYmU0
JXQblKkURJ6mKC20YUVA41pfdsqcoIAR/R+5D0a3lji0eiG8nGUyG1Fs6VEBcIUj
Bb3XlxJfd7hY1L3JGBCecI5Ttdw9W7EvKa3FNd65xstPdqiLOotas3GNcpnkpxii
3/bpzZNJO+YPW+3SQwCvIIH7Pr9+Sb8UkQvyO3dhcyDBgvb31oQuCc9utCb39ohO
kCMiBRZCmnxirMktG4ZtKNqW15ZhJriSNsOBnekl+65KyW7IS4vO7JiQAbAA4xxM
ddQpLVo4Hiivj6KEAWY/AwcI8auaRlDm7QyeT6Y+TojnJ+kYDK+AUGRq/S8R8Epo
ZK2vaXdTN0ULuD3umBI68Ihn2icPUzOgM4T6pfzfnGfM5DMTREEzq8CUwrYOgILl
e9BN8I+i8WJiw3l8r5RvYpDTKQYhtIc/UoTctRKavTddRbHaO3K9qpHyKBSm3w6H
no/ACLVOx2mxpDTcpWJcuYQGQogIYLFvQ9ETBJVM4sr+WLT/G91VRLb3hAPkyJWJ
+5KP6avA++qShuUpdXvT3NOX5Tb2XhF2vIKNKWHt7Ccwj80SaditM4uxQEWegqFh
7sxnQSaOqdA1ief+JklJQ8QpFWaUvM1QZrRrqIoNw0Dqr8AxA22FXVNR5DZowbYs
rkXezcS8Lgi4KquKZyo62dzWqwe65FDwo/TCMZOOtn9r81cnFm80Ka/n66QFPtF3
EXvOy8sklQwyy6Il8z88mJGvVQNMmuqGLhLKQpM8rkHTpXxFd1zLC8TihjOQ4LhJ
iWwsLscUYnTksBM+1sstw0qpAC4jt+t5EpOIOx4SwQ44ALcbhoU4qSO5Cl0wrbCL
6aq9kICsmiQMa585WdCjLUdJVY1dXusGfr1Q6hPIeItAZiAUZhoQCOuW6MLPz+bk
5yQ34hmOijhUzIHiZ/wmgqmXwkOLiQ4Zj9QAzvWAvm8aQynrB8IZgNhqMIQSYg8o
GOx1G5lk8JURZ93jvUntKiNsDeLWzVAXVjAUSe0ZO0ekzUUR2Tnf5dIhas3XSG65
8vTcC2M+N4PthX0/UNa7umAtZpY8/4fFPQVDgV7fz+RLKSmJwmJdpJxhFtiJN4bR
mUHswLYB6jmpucakJIGEyoRYUa4DorrEDSZkhcm82nhkyKQAEhM81CKMD1/0W11b
6zK96or65kVn/313GfnxGw9liEkd4UXhT7VI8LD728OyjjpimEGzpDPl2skFckUQ
NIPFy4WyQ52KlwlomYQ7iZq4gcMX6E5GWUwnNUSEQmw+w5IitLoWH+Yqm1YnmeeL
0sqAtO4ef1F6jpcdkMDsvxUG+d+0Jv4EM10sRZKPHH1/PExaH0Q51FskZAr+AEO+
X34qUsuxJQk1tuURJ8cqE2OXsaGr1fyRLzbZfeWOx3gEjAgO6uV6tcdeG46fVCOe
jWPa+8bjtwIxjFYtWHE4ZzB+2aVzJmWvfD4T6ATFBOabt1+Uttt55fLsoKvJ/33v
vqeB7Oy8Q3LKBfp88sQ8yp5rVClanIoKYQdoF0F5aTCIGrDRTedPiNpWurK5+S/T
+M4SmmhcyqKumEkEi720nyCq0qSlL8NVHkIDibDjb0MJqr7vvhX30Zs81eBioA8q
cYEG9kvdVc2/uQwRUyOVWQxO81icx8JplC2l6o6q4WP4QJzSTRQluOXlzP0139hs
+pZKUEtK8p60bS/DxyUmZNE0WgYKpcEuJpVeGHCGYMIfHmKYKCiCZFly4MrqdruY
oImX8WjlVpHjYqWFGxjUPyGi8ramDvTURVr7+FQEqe2Us9uO8sqfTiGinHCTVJEq
kGxRcNwgipbtr7UZ8iGHGtu/gbW5SDexF0pzpcEshMiU26KGMGFROYtIDgweigP6
74zUr7aqe6wZJcPZiSWhs3kwcDxZyCyVzUZhX5FTUUc=
`pragma protect end_protected
