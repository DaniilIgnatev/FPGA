-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BZyHRC6hfFJtvlAumKdB5Xb84uLmNOAIV0Wx/DAbcEgHO87FyI1fTui/kjCuCyWAJQdZgsQvqRKF
2hVOzTaUxrMeB6l4Qyr7Z1xps+6/VGiOCC75VqJ/WJZ15v7wfGWkPOZo1wPBXg5Pl88xJj0Z48Wx
Pjc2xGxbbCavtEnDNsftCslQnohDRH2tr68u477KAcQYhxNs4JRgPjaiphZp1NT9+D2RYFQ7+PJf
jklC2p3sVNAQ3Z4a6B1qwiHF0piZXUH01pz14k4a5ZD082vFXoUH4dN0kpJascd0ZeKGgDc0XINE
mZLcpZoSBhylEu1ZKui0mh0J+3e+PyhYk3AAdQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7296)
`protect data_block
RCC7NlUr6lOoQaM+tRqBT4RH92O3HC3zlPOPaZdHpBJ7NVV9cwlW0XBqxYwpoTiZE0sdmpovCtLf
uYjhYcqVgY7q09v05xHA07BN3OXxUdKaDvDhmPC94quBu2O4KzNSbPgDsxBqWzwbX+wE99l7EFIw
J9iGJbcuNoIfol/XEea6WnDBsiZNFv0GUQecVILb6GkeUol5n0zg2lvwzyzPohqHOx66l0xT7DWd
Glqqlzav4rlcLaB9bBLWW879buq0sKaS+ovJKexaCPwOOTTi7LDsY6sHooY4ozmx7+i7/rUfbXKb
c+rvKOYfnWnjqmG+jzzZKLK/BaSdF3SmNWEruMd19DM3+rnSKpCWJ9Bs1C78++/U8u/AyKgVWqdv
1mSSrAnxeik9PtKIFU6mjwzMtl0BaWTQ2fbTWqOzsDTucBMwGOZnMLlFXzW4gkiS80wxylVRVi+K
+X+hjt52aBGrGVolERiaYVf7qUjKDBCtWxBWu+xbVDUokuUjZIkrkOcl+WOgcc5ZuAosYXWHNEnF
olHjaeSYTYcikMDvniIG5iDOLjSlmPBc+yXparI7yY87pK2bcxkcL8ve0N9GZ622EkOHlYps973f
KN1p7YmvqOBQpx/QjvCd3bEnYCtPr5wvK4pjyQ2bxkehvjPrOGe4XljELPkhHomgvHf1835JS8RJ
qjfFAFAG4Acx4m++N8QBc76IgoX5J1QesPSPWY/Wv6YwGPL4qqdj5nyWEfY3XnRb+2DIMzpAPREV
9qftm6OU86uIBegLYaCjT/0y0o1WOQ/7d1qeyXEQOm3bhyrFaXsarcnoTlxVj2Gq9vQ6SlFk/0iO
AV+s6GlN4+V0HzzNv/MeYCukxqfAvJHnImFJ2E3peyW8v/1qpXo5PzJFtstrv9UdLbmDM6/M7re4
dPb0Abk8m1kJxUIO3VIsAGFfgHjuhaA2FAwuE4wOKmDzcIpx2TpzI6l2Ske/8WsNFna1B3BqldoT
RMWneJ4UmZZnrJGBtwq9w7E3eWjK9zzvYg48NmlByaG1n0/gtX2FFMfLcUfVe8A2v5cpaFqBmL1O
CVn0oS1+Pz23j50w7iBUxzbj4dm1VoE1RH3gMLceFypdcZWvR1DU6qB2ImPK7e90/YiOfhYHEqBf
2hRhHMaKr8rXo49uwBRqdt7fpWPj9sMntzunvehIQSFNKXvZourP6CUaS6X/7IhUkr5EGkQ3LcSJ
LLNb6UL0+nrnDDHPJZnz/YtSmPg5Z3WTX90SuZ3+z3mKvZAt4ypZH3lWv7tmPM/YjEFcnnj6o5vf
8S+CAvyQfiuv9aygzGvNTIqSARhAxePF611e3cQmiVE8XpiCtE2P7c6Yy9yl1hQmD79dwP8BT0EG
Vp907D08eJvD77I5g1AbVGwzZMCfQKat91pIDggcD4YNEy2+/EqsqBPSfLzwRAsx7Sg0zhzKdnZ0
duXFNSPgW4mmDysGOWhA+IAeMAcmrSoNefm8gJ9fbDpBqFe0ThHIdloCAjR+42c9+BB8rJg5Z4aD
GrDpNL9782gC8B7xM3TCa1ma5UFpqxRYasoir4LNWL0DFe/u/87wMPqaARFiDuaU93LvPJ97sp0d
LHKnb1hydqRQzpZl+2k/iU10RhSAviP9M+nof0mfDvGrKuqpxSVkJwIG5irPHo2R9JWfC97yy/Cz
eCYv7u5mGwGMqhoKQD5JZn9gHfEBQ78YlUW7S+Sk2aJbXN9sKRR04es5p18JinBE7vwBe2O/MkUq
V+w0DUjzaaPN3L2LYuB5yEOSF0DuQfwQvXB+eCBIQNdw4dbvvMzwIdoWvEwv+0g//awvoDFDYDd9
SCCJPc2rPgNWcokQNDwUtB18IAbU/x/BKTIo2/QtFF2Te8L9+hMTYR5Jk3oN5IeAeeG/DmEJRrVB
q3Zg852c1/WV1w0HAgPKgJuAXSNyz9itVSuVoUAj9xTMMyQ9c/UkmNf0/gQJp3dzNc1QK4CmMUCH
QEdWHycEvx2yMrZ5AJsU3vr+uxudK+TwtmicIV3oqim8hBSLaYWErbqtL3lKilD/GR1l9oSeqByp
fYAPrxqtmvNWQFpozX5kB5wIVhcd7MJNlSJkeHfvFVd/ROb117x384EP+ApBjcu3yBv+7UfXaTKu
um3Ya7NKJmzOe9HOGfDsH2IPAc5ZRcXl3ofZ3c8Grom+xVZIF6irgWj8D/O0XetGHezR/7gg9wr/
qvLk7VquERgcyciZLB+1E6suDyV3YAE7kQ5VhO8BgQF1Er0vZivDG2NxcpgkT9vjxUSfFB+waEGS
LcngrV9ZrD6dwp4DdDmEhw9Ql6/cyX53785zcr5aTQ1dEG8HZO2LGBDHboam1oxS8IDvN32i05Jy
rec/uUQGf5Znn0DcVNwqkZzty/Yp0q1xPWolL/PeiLkDeqXTsGayILq2YLsnbTq0bBjmJH0TR/lB
d68RxjtGhbih5LcJ+C3R0q6YeLGe3eACPmhfk8Pv5YiTdm2H9K/oxbSbkZQ8wlfWmZDhno9nPDuJ
AraiSqLFIXZtM2wRWjv+/+32Km/gwPGPrJaNyGBhKmx0PBVJpcV9tbF5Af3GTjSEZ80NKJ69v9gL
4SJKAdTbk7XDIeNs/lu86W0dl5tcQg4BbfKxNSu00f6RdWUW1DTTLY/waVr850l/mDroRABXfgm/
COOFfewISd4Dpx5oEamDZ1GCPrr5xOSuSgtJAMO2DkNHnpt1dU+GD5g/NR/6Q93H3g6H8wd196BP
C75vL7epYNT+0tLFQ8c3V2WUqsFR9MhxHADc9uuTUN9qXrj2owJuLOF9AC1PhtVxwaSRxlUCNPk8
dyWbeycCYl1olwA2Zoh49kd8/x7mY5GdvTNKGNbc04A3PtxsaI8IOLAdyQvoqXtK4NyaVmhY/Ak+
MymBLMC9o+fu15Nq6Sps6jH5DgkSO5/2UzsZeqNrWm8pn5LGbYEmRyBeND3ODWTf9T7wQdt0z0f7
2T+TEF32LxvKH/aH+sqhvwkUfOUcuaLty0SVm3oi44lk8GeciMOh3X+p0PJ0wNYBOU5GIqAKz19o
aSISaQIV/8yevT3RQvKAOwqinMmNaxPGZvoyaApN/p8arBN6JT82fXCvTMZosK+YR5KGWZwVPAq2
HDCmA76kv+MoGHeczJMAmlK2F++IqJ8OJA5xoM6yy7/ekFSo8i+P445K+53c+tDSi9ZJK8Uiy4Ed
CwsnuTeuU2YKZ5gP/54EuaQSa3Z+fRDnlLpQmeH5k7eM8fQ8mvPGwxt62RqYqP73JFHgACUceL/I
y8l0p6go4kHDy05kIYRD5kkbZw1bD+uWJJ9llclm9t+nDFCYU630RuS7/EhGRKo8mfaOcuHF/bTJ
dQLzIicW7xNBVuLkbxRoKdDiOZd+a/vt82IoMjiSoLtRwCuzeEhNZxXdljuIg4vK5gkgQw6soA+H
VtSQuA01JZihHMbfrvlXCFVcDjXv/RlNPlAhqIm9VLRfFN60iWieH3Un71MNNq0glwjD8T/Pdord
85d4BP0zT0CGsv36c6z3tSePkWHXGx2JyrEXGRhuDGELiT+oYhdmRjVs5ZNm/Wdt6WcM2hqQd8NF
bmtXdcIDP8fh1jffDT/Be+Vejf8vSA29DiMmkKUOvDjdWA5OSlvEc7sDyUawn0e+yHV0WsxdhTFq
kQdJBOzk+Y24A1NEn6Kgtnr7Xxsf0I1Djrg5SbYEaM0apHU+YMHN7NtLqRBDB4iMePDwCoXrpuKM
iKE9wGzDnflkjQkB7efz8tFVCmYmux11+FPMWX+uMH3Jng5kVTBwkzY1qbieExWiypR829Jys0v0
NLL795tB+nIPDH+Ocx9+buwgplHqQ+/I5TBGi4XQFkNErj/MNF295X5PnF8Jqo1dIpUAN63BUXlU
caBSlaZ63mEFKWh1tG/Y7NUATYFivGAk6z9LKOi7o+0Ae3P2pozDrN/2lt66HOmaykfg/9FI25G2
+t5G1qGMi0ES1mC21cAz1nnHj2gdewytPb+G4OfG675/as9qMunq4Lkcg6TcqpKwPqAbXMpm4pGm
uAXUo2jc57CJywBsp6MaxWruOiPDW/lQfKG6M1PZp+aNRovW6zgmqRYFf13KmNcvjA/mNrrCFIx3
CqhsQ4OdcPuXfecdlYU8xA6FkDfEqfDwMWwBTshjezjaVYfjairAAxJEv75UAkbUvhrSB/egWHhr
j5WQ/0pBsIlk4Hldb/l0NKppWnbObwBhm6wGEGcnm578lmdGLfgEY1IZ7OmtqUutMnxvAzICf+TQ
5x6n92G5gSq0Ip8mclkdOjGzJsGQi0nsvotHQVg6GlyvGaOIZ6FpqL6rsr5gwSfMxbqyHflw+/P7
6cDJFHrAIB6SLOrjbvGJEMNWu7m27GbNAI44+hUBRKBSoBZgffDYNi3a+MFhO/cdI3OET7oKrV1l
uE6GX2mO8iAnRDDyIO4+JIJ7OEX512ioG+bhWXqF2JNNEORDH+LYIh3Lh1Ywaf0hufgIEEv0+Hh1
jxMtYE1YBR0O/nizlU9xXI8iNJDIhf97Wz5exABH/ljcQj5VHHlDSnrgVwVbdvGVIs4iJSZ4HDct
bIT3NpnTm3qEoLcfJ78UeJvPQQF9iPbnYLzo3JmFYdl9rSPghQpIYn2pJPtabXQt8OA3Ltb8txPe
G7wi0+ES7eYCmU4DyzL9oV+QoxKIEJL3qM+dXT/0nSiIvmL4ynQwC2BjM/N35rCU6arRixwyIE/w
OYzhm5mMP7qIv/abxS0ul+FVPUOIjhY0ra5G5bi35UzR3dGDTEbLaIZTHDJ3xd3fUzdxmYa4sCmn
ruP5AS1kpwZjFZD1FwdW+HdH3cHoghWRy1IjArAG7YKqK9TCaNrOv0jKENBt1K/pUsvDbl3cbhvW
6GgKFRpHkCrshtOeQUABejPp03Vtv3NQFv54XAyvMNmZqOpYqT1HnI6RN5frQX4yFUvNubl1j7aA
3gZFezcwkZevQmPtqlH1uNwcScNkh8R6CGU8St8GztcaZeipAXFSO/O01BGknGc+11pyJly7jAxI
ECN3A0fRITCQsHjy/ADTTUNCjc0eEq1u9QoJimwNpGE20o3kxJSN/K0UZosblWACBqyJ/AoA6VmD
/M8c0gGs8pieBbuFBwxbv1lhAgQYQha9WTL9Y0C0XOApfPRnY1Bx4Pr4Fk99JH3/0029AokPB4Zq
+cmdr5dizc8JM1DikMnnLG7/iccfrDr/2JkFQE0ZYnNSPMH2NB/o0A2SGOYetrkLbDqRfgtB81aI
Apww/s+tCUNVGkGQzJvcTtwKERmnnSLeQOVVyGDMzDEvntjzcbOOi9UVmtCTM9IjnY+3XBTQAUed
dlvJNOZj9g2jEBpwEQmyt2xGoNtErWeEG0xMkwitCpaHKXSZQ/VuA2N4AG5Fd6kGdSo4mF1D84U+
1EqKeHdkBvZoQRdaqCNXBMmQchIfjCTyLWUPwzpqNCNo5qhjMfQOJA0heGfciMOcnHHan2zw3NFT
714fP6bYUNWE+Oa2xS9Wzk8lufuUAknxpTQ8UqjV62u5dSZQ4qnJd5PbFo/W60GPqdENS19Vm7Ir
qEDR5uVYvpKAkG0Toi9MdFqo2OdMJ3kjncnQlPnnaxeKylTAhQPi6pfC61FVv/yez/Qxf699bPqa
FEFHsJ37rCCDSyz3sFJEBRwPYpjk8XdcX9+8U56Uy/IiPMAl9cssT7tCLuAV/+Ldxxe2/kmL4+61
NMtlIp/AaNKmP+UNPFvEuoV//K67K1vUIdIUZzdNMOuZbiCJ53FA1G+SoOaAONjTW+K/GOkOsoRY
hqaxEHiFdmLiwLmS6GebFyRPGEc4knEArJA/U5ZEIQWdyA9J7xqcJAXquIFpP44Vw77sRUGIrKW3
QfwmOr1Hq9Rfa3749IUh/P+7nTC03fsXzir9w3XF5u+dTdaEbuLZMXLtOGlgp5++/l+OvDcSm6hs
Tpq5FNOhifARub4lTb/ZI8EOaSOQkOVE1T5ToFC6NS0cqZqlHLlfuLNCEa5qZV3MHLj5fHMrbO5V
4sY4D2fmgBgfX2zP6oGHQdEh94V8xYJpKIOzqOL12nFUWCur8XiWGN6E6iy/AOCbSfvsdRGw7kL6
hoODSkGqg6V6p42LZIOUA7PY8piHPoTgjiUSFTEVIJsBarKdroS4W9rmuZ/DJQ81H29CN57TpoWg
fM5X5Kv4y1GdU+a3L/cWHXw5NiT2stD/P5CQ7GFkhegbfH0uPtCvhmK4IIVqzNT+djJx2rxjfGVQ
1F0laFF89wt05hP0b4IqBLTJpmgLmSG3X6aUQGx6BgvWZfB+6DgAPq93TUG4ntwPP0SVpPdj7m9+
j6uqkfVphRyIwH1pasi0q7/E7IPcYqlh2Y7Jm2oHir0/pbfhoYyuwlU9jqsizm/ssH/3F7Ohu4PZ
0e0/7A07OqLDFG/52Vg6NXPxePmhEOQRfV6h5TT0YvM4+NqPelKB3ZX8PjO5V3223xMPqQDVQFIW
CDrqSLMTn8cQWMmocwLdCIqd89G3/3830AGB8b6JXLNEEbtmwPwAOGABEjYSG6WFEXRtsa/VQ3Ba
xuN4fyIr8eOCjXAEuZH9fN3DF8j8JAiike9O2d1vgsTxhASq5PxFZtl/xFTW56aDmAM8A7MnhpsP
VEHybeCDW660XlXbq8r/QqHFzzTJBq+tnycrh2mTc6+cmc3Kaf324LWcJYNCSnvdzurSzmZrpysJ
MrIxlDTLRGjKSVMXwjKnvOWqsz7RE7oS7S8dDyX61wKi1+6dP+NVUZQYDP8h51xD7xRdR83BDIT9
/e45j7lKgYksRdBch/4VNHSL6zrULNQpcn3BBgZNB+yPoZe+Ej58eRAzzHB/SlnG5s3aJtIwbIWm
KaeBWcwnavH3S3nRVd1M+79Rjfyqaw0qXfArzIv0Rz59yyFsWTzfUw75oa3DtPDk0qAE4IRs+C1t
hg/pHruUbL3RJBb6e0i+O7mHfc8COHalTpoA9bA3cc7gtDqI/2wLaeftRTCOxY+F3uX+i3pWR1WM
/Svz7eezzOvfArEzk2u8RJcC4GqGX9p7Z5UOFzyCJLnRpXsUbEpj9l9Ts2/pvEzknUccy+3G5DmO
v0Wah4xYAn0Y6CuW9t8Txp2Ijoi/kxRBSllnNDvZo31aqYOzNROUeSpNoxdYJ8GywZ6h3/Z9qkvw
BM6I+ioIWS4+L8P3UA2kIl58mBIR9i5qyo9xOsyBqP7FSmlht35rdQZe/abS/+5D0/yfYALVG+iN
Cc+d566iJCrcY7DiLGlC5gKj4YI8Z33CxdJnKhvmPgJPYUbRo+HWKeMkxy8LdzjYH8pn0jokZwbm
DXnwZ9q2m3bIUWQpgK3l+F9+one+eC3PfFoYwBYqfx20E9PLITm8VtBLFsn6E32H0tSPPb8RJs5y
HG8hemWI1/mYPNQvJE8kS5v1nro2I1oQazShPBHbm10vDr8b7eyb8EqrBMD99JHnhSbiuDcoaVE0
7U6a52BVNWCd0Zw+eCNoL/f4qUX+U7l776jrwJ11+dbVd8oZLQxNi4e++1QuXDACo+bdGK+NDe4p
EUIHj56biRBeg8lrPzxtElRHrH7oGrf3vsTqN35pThIeWCm7huF95q+0NfNvw7IzKucmIZtC+x+S
nwBuMMag66EWa8JYlCyo7VWYspPYCZGTiDumHB/NS9tf1jVR8GRF2L34mjAaoYm800aWmh4Q/GHH
eoUkGyXDWJPu2f4B+YvF+jk3q3XyhtYRiypSrU/uWTc1s3Oy8t49bd4x0fEHDFu0tuC37Z42lDUF
XadiE3WItPQb4gofsIpbO1XYWd4Ap8+gMfk9vMQh0D5FbMAO9fEKufOqbaAnUXJBsT8Vfpm4ToNx
wlOUijnq0hfh3DcMXOJss3zNsjBOjjwznmqwE/pIgmtV3aWS6lvOnUGgr4ApwrejmVBecou0wcL+
No7+0f0tF4WOmzPULnvUwtw8X6b3lv54A1J1Qh5DkuIIYJ82iMD1G5CKRdJBY6Luw2GQ8596EYnc
K9Fc7Z5eFwXLlW4mXDaUTmq2USiI1dxTVF59IWlPwqu94HNDfywxGJyS9Dr1jYimJd55bnu4X+jQ
Z03EZe/AYdTMepQmoAJ9uabKWdHSWfCetZEroX8CrDEOoKQF0sMjoXzCriR/RwwisBnrgfBFOYJ9
K6A5nJXxwRXr4XP0mvqNKaHxrIaN+G1UKsc24EMS3/wxoj9m82myPSjvhrHZQQI9Wa7oRq8GNA2r
tKq58Wbd3pE2o6bapNZjDmDBgwnCaKLNPN7NKUxcO5Ddf6at6A/IB4CTlg5sHVgAiSeQDo6GcqOE
FzyM7yA7vTqyNde1xPT1T8ivoX/H/hU/pIUS6kgINjRNZ1DmEp9ptraGAuZs6CFxnP5g9pTA6B8d
mDVJGMP9f0zjKH3w6v8v+QbWcaWDJrc554wOLdx11vJOBFWl/e+q8NLmrJ2kGjNW1OuzRqTKlSF9
WGi0kCPv7Yazzz+SstGw5cr9u3QBhNPkvt1yo998yl5+II5ipmjaptdJ8zVbnM30ngdo0m+OUr+L
Y/5j99+33DLmKBK2J48nNF/E1ccBGVA/o7vLH0zaKyERPFf+NWuk6SepTSaoFe9T5768PzA4eJq7
CZIHJou4muX2wTkOOQ5XV6j1n8vT19dXY8YOeeFBEHM97b7iPY3lWhXqpPPdO4eBtFsm1rJDmwaW
mWH6eyhIbkvC0TGJkV1kcJbD+bJCh1fh/7AA0rYn223JSNYCEe/duHn6VidSPK7S7ZuwlQUkV/Ks
PcDiSBSN9gyZCuSpVsC0+JZVa7QtNoss8QT0n3u78y7gcDIunopXxEkMZFuHPxHPzlMgAjXVq3fg
c2T4C8c/t9o4Omhx4lX8+gkEUMakF+ouvaY8W8a0FNH92vRfPj3RoTHaZUHFk8EDJ+P7nb7qBoOz
MQ8o5yKhhBo2KpEEOd+tM4gzTxEUw8ulWt/8Dm2PLLeDyoFYbP1FSdw/xu8Kw8xAtu3kC8Jm9vt4
hZhGXXc3tlbeqPLIwREU5ul9O+oOPCVNswcvewvfi5s9Ebeyi8VFmyRc3vbZH4nbEaO5JKeg1YFH
LNfqt5RuPrUvz6ge4FsEqd6pb9Wzts4g99PfHvBnLBT6kHP2SLUW85d+/E5Wzh0rYgwiD3i/96vm
Hv1zBiXdCc5JshX6jt7PhjmchyrTvHHD/tGCcmivJwZqkFaVKTQiO2etwL1GRL7kpuRn/i83vJeR
SxHHwO7Qs9KX+WHITPDsv8ON61VE+uk5NA1SZDnxgOZfduRWvQMsR7AdNNuIM3lcHb3DthwGutmM
8ZEYCNvwwYFqQLO3f0Q8PkYUwoAKiBH1JKkGkqU62nmW1IHohf+oHCaPq+fPyY9sVbh30M8kqaNK
zUnqe8kKl524T1VasJTTOwFiD0d6iaEOMi+kGmqz0+IW8CnYtfAJtS5Cz8s+QK4wL+vqexpF5gww
hKaEZxhPauiKl18ZmMxjcwkxBeIhFiVOAW2KYQtEt1jsjiBkjYFYOP8Wv3CZ5tafKK97Pu3yqFWu
euzHiddRyrvcQ4jmR/yVDijVIFD6qR6iDvaGlnodcX51onTPr2hf/aK/mIR81TC2pyXEZPfL55gL
ydI2/FrmoJcvFaxs53rmxWcasgSnCgyiE8A7qCTixAIFr+8ynwj5Cd16L+QcuboDzMXU92LYfIsr
IHDJ7sTgolpvllT6rq9rJSMf+eZBUEu7w2RTOwVQ4h8M8O6vq8kkUO4yodFmSY/dmS1b5FHlUkN1
`protect end_protected
