// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Tem+Beh1RlazrfWxIO4baeOcI0S/Uf5Q7cMojCUZVJLJt1BtztDkBCvl35qScmi0XCGD0kuNmY6Q
Ix/MqNFm0H/Oment7qGe375g0jZUsAe++4SNz2yUoAgDsfL6ukGNEl9cjTCoi944o+E1+SzPjvfE
m3AlOwVLomw90H0PZdYtxYwWUTNtISVH+jmhFobZf5aRQjGVt+DFoZ49Yglf30A9FjdGU+XtWfp8
y//Dr8IoSlcUvV5vGPystbMu1ezokl0S7qF0n8bx4HFywRQllTy5NpRRIa+2XJcoY6M1rUxRuD0K
zsF0RQDci3hS5Nz31RvWaYHk/702aRDsbh37cg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 24432)
2yIOoYPtigfmfxIjOlhpNu/IEwen+T8XPsD49ejxhh15avmARBwvcjHh7FpaHGbQnlWwkmiigZP9
VDTR9S7YCDQdageJQ3SWPl31XMsmSc6AmbyQAmJRYHP6dAZ5u1ZdkrVHConur38v23xxt8FD4efr
T1sqVDOkugFLprJMQWPzEaUyze1jVW+8BlTgAO/O+MU4tTb4ruXDd5+i8rfu0i8UWPCq1GOgwc1y
TDdzrIpkDgSe23hKDZwXvuyZwa/ydaGf5zLmKG+qb3XtKWgIe2k1mJ4jsFzZdpFO0m0L5jjukEpk
BVgScLv9qtHPxOtIBs+AsAGEvGMFG+i+bVyq6yB7UvwbV8JFY8R9VhEu//sfq2j0b7D7/P1CXuP7
Z30UpJXjpt7Ju5phBhZnIuT3o8+5RW19eGC9pSfCDoG8oLBIL6LodaGXUT1kOgHqdLYlYmkD1H32
6RAzR/wSaXGEpJKuZfzpbAd2w48YdGsYZim5SGg/D0PAxDLcl0OuDqVwlxBxWnwOltVcDigJgf+O
mJnYU/vHL1pHGIv4t4lHUbfpKLfYUFEAw0XQMwLf1lg07EoeTgfjhsICdScaaP9hcZaFLfKHG0r/
VunCM77MXr4ycOKdMM6TxE8LQJVIb8CuwlvgUcBFm6rqpNeMnom4LLmxMi8SOMxgTQW0fWpUJb90
4n1H0P/PQBraoj9iDs6kpaF7pfHh7V3rNhQinmKiHTwakEpnezLR+CEaRqsJ6TBBuF3ftdU7d8lu
4G5eDfhaPz+wl1TGGA3VwFB2p+B6OBauVaji9amLzppmPnh4LTaoDMwD93dN+VWDaRkeACsMYYqn
9j0CYuv3ZNQHoRB/4WTyBQCY6T4EPtNjX7OpWTaow5AoGzG9lEG4CECHLdR5dEid1d3427Zfnfr5
0PaxEcxRxgX69mRopV9zz2/59wJ4BGm69rmkpV3jy/cIDo2tX/6n7LWfyJ0mt+rDL/lPThdk5St8
EyXQuisY5CbIOf1zqZf/L0gZeat5Y/Fg03L+0R9Xwq9dmuHprKjru4AyNbUqejHd5X14mjcfb2AY
Jf1lNnEUVrB51Krr7Z4Y64PayA0zuhtPFj7hMywjuaVab8y+37SWpAcIsy/14MMcG8bI8s6jnDlM
WM54+tvqZzFGf8up11EFTi3GWiiIbpjAzeS9mCLNSZU7Gi895Wlvoo9yQmE3W7Ea6PJxIn55J27l
BocZZWbrBjTCeQFCDT2sGJblgomqkQOOyMydhf0iPzj/oJUqNERYrxdo95tdi3NGB6jkuc9+lODQ
VBOJhjJzJruthPDXFUP5/zuYTLKPUu70x6WZbMc8MSrkhlhUCHm0uQKnHLgL/B5n8S43wKm3N7xU
4g3n+YIp7YWayIQ9yoZAvZQbwPcSYM4LrXmDfRKpjUYc/CdzLG879r2H57uiAvKLfZTwNTpAkHF0
IKzGqzFiAXE+U8wLPRDSyKEmHa2RpB2JDRKD5TsTbPOjFGA6zOXo2rTKGQM0XmDOEt5noX9K4Nyz
uPNYCQKikuyw8btACeReT5I4VXmw0JrtUr3Fk7Lu6abxLjI74I3w8tjcoDF/Elrm21iKj0OvlFjd
SIj5XWZI7JUmY3Mg77ZFj9fUicX34zjrxpAMFxZgy9YQAMA93kdOhDnpbHYQGqihAZGlD1UnKud6
sK/YqN4Q0KSsCJ5xIVx2eW/IUYRXbl6EpnCkm6gf1agCYjiJ0sMTIh81ysU+PzlcIxCTU+bJz+be
4+X7eRNkciFlRyyzgTBMMI1Do+G31NQEwCKN1bKVCKdez7kl4hr5dBE7vCoiVhNKkEEaenZb7HmC
c4zwv6OydwUsRi02dynldkn9W4OlZil2h6KwLO5dYntcKLVMvdMSMULFIYjCcI/5BUm43iORkcV/
n4216RVkp5bbB3C0cMnMfOsUjkcnyXFmyUnXF/SOBZLaNnOzzZzHQ81NKmkZwvK7MeD6mABd3KbX
nBkXO3DAk/rjoRZSOJsFNX14Lk8U73FZBZTtri836uPSOy5ZGGroykI996AFmvzNrvoMeBLEKOzC
lyJ/JfrY73H3B04ulpnFbhpX3qsGJQAuRgWbGuZ+rx94zi6M2kDnusWP2y5X1cwEr3pBx8GXzmiI
fSj7a+23KN/8c8P3JbGHGp/2PZJUAOSunJ4oB+AYqnUP/PKRtbVT0HqOv6jKDYxaH+gyhfwTOzK3
GzDvu6XNlYdLnWgN4LVoDdmQekN/8NO9WpP753o6nYcHoZae/S54qU91eib4xO7zYIXmLQXbE0iJ
PzDFbWTIOHFf8mWx9NFvxNskCA3fEpqUwzHLk9wb9ikubenKgo7667eHPTD7+jqu1V7ZwmoLV0j2
m4T7FEUNFE685S4Lj4NPkMufroCylus0PKlVmBHQEKL5NhbnpbyIsW9ZeNZAgtgRVQALTZi/ggPB
neQu8X9/IbATU8d1+VuTtgfSnM2ecxi25N7YadlqgUp2ENOsz+YY6u1Vg2IUldivW7Xbi9FAe1f/
mq3ttcBISRW79AhykbKDBK7gcZei1dWqRz+87z1I68IUgF6qGdaRg15mgIlHLc4h89cTj9zQeTIj
+FFYi16+IQevajkxU98q5iHN2/egPBE1PsRUZbTi9oTwUZdUoGRM3ef6xCHoaziVWSCfrmcL9sl5
i+cvkvXrAJPtzF63/O7p5Iqdyqt/qLAXTs5sOgkUTJmDPX/YPsMKs2yFMOsCDTfvJYIYSsP3Cf2o
r6aomhZ8lR76Jyi79wWm9ecw/4lLSGf+PEfMGvtNiKtdwisNNafkUcO78f/HhYGuFZ82uVZAh6hl
zcZIHZdCMylnhLYOzGtvgkatjdv4We+4NqldmGjLm3DPCLgE9u9349s0ZE0JfIlOyixicX1dg2LI
k0tIR9OGgOIcK1P8dxUySF2A3z5OXfdm5Vzz0xjqDa3sD0ROmUsaxWm6YHRx0+vfUfmWrxy3ga6V
Q7xMJY66Xf6RY9Jstmb5I2PrvsmwFnwsCZbmFk7+dBpcOeIk9egzm6b6woM345uodmLZyDEDx6FN
VFQ2GiuTNf3bKbL49ctWnsHNYmiKV8P+zB8iFE7GWwjXhGVIKl5CQc7zdI1kct7cR+laC0XgqH1c
EkNHlFoER5DouGua2zbYss46vrBcOYQw+syU8R/TGjLknZBgXUNMuyg8ReHnvvWtdfwbwpGqKtnX
9ztlCo0F/KgGD7yh4tArkAQ7MzlWgyMZg9zUKtW8Z0uraRrgUGEBFT/GNTs7c5bgbi8n0b3I6Iqv
6UO8N2MtPVLpuNlIlHrjecHKKaMopg57244Ch8uuMVmAJIJOugErVOheSjdWnIFyzliEVJY2Prjt
ABnlueoS+h3EoA6tyIK5lK3bKpi9U10SAtZQZ6tAbUElA+kbE0BcZMNe5magmcldzGpfYyXBto7o
A+P8J9j9s8pUPAF6R27cw0QX9pkdCcftOfPWyOPpdtTIvc0p6cNn84BNwvnRRhVFKQxxn5gj8bH0
qVWZlyxqKV03XOEY2v0IQ54f14Y3F7NVTDwQgbSBBK44tz1s2GllPgwsQ33eV8SwVauRXcw9dOXi
H800Nj0+xktn8G/VMxyFjP/FDD2pSLK52XJj812VX28IN2MHCXJPcZBDH1Ha94xaRLFCX8gaoQgh
4T+pPE6kvIZBe578lpfjFuo2qk6av2b3BAGIBUASzy8dLSBgQII5nXJDOFfDFpag9Fr5ov44AuKN
+aZVG9CQpIIo3GUC1xAz7qgmU/L8XRISXsPRxLiZuL9P6pRvnRcyaXhGRAh8d/ggNvN8h/5t9Q8b
A/eyLKxUMKOEo7nP6qlN5yvo/Y6wXQFnVaksCCEOjuGegDM+nWuXxHWnVDOIGDtH0xWrJ4WO5pqh
ECNKobSeg4NrIruNvW1TuszuUaSQRdQlJJ2quWh8WfNHquUqGSGqC0wY3UItNt6LY3OeODKLGn4O
lLjK0AwOphdKS8rT0pbAXFrtKI6hzlnmbcNYjKtlxyQrylWAC5lxX4tFDwPv0mNRjCmJIwA94QSd
4kSPMrMBUs8AaC2/kwHWsge9NzfYa0Kqa4+DlbPo3nUPlCLwdqkcljhfnhpYPvQ00b8Cv6Bf73TI
V0ro9kqV6yU2C33qMNaf4ur4MBNIYUpbow9adnRll7vvi5Oj7fEt7ZaRHArH2t/f4zyVvq1pRffZ
RWRe6DCzZbJ37l5xoHCDowaIWJ574JosEURnlPlF578QhYOHDIw9QB5m6LuMZiFENpm8QlkwOERA
0Bk9Y3Qw4XKpLNhDFomXq4t1UXN102EFs1T5hKWb2BsoHGOLPWyiEnNPF4HG6blvX0HOrIXwPOnz
kswpseMY4iZtDUL6bBggtVpcEf4sC66ZgWVfnzLDuTeoXbUdOsL6z3PtVBdIVzEzPzqdo3EdPvRa
PojemD/w8ikEEcF1UAqWOoW7J/zF3rfxhAxFZDD16MMLRKTOTWZ40tNatOO4MrPjy1dn1lol/ZlJ
1rhTvABYPoPQ7vJs1Fbc4xppvBq7cbbLiAMqx+M2xzPk8JZGCDAGhUIVwtbARdBiJLO+OGQtJhB7
En2Ah6Yg6CAyioQSgzxEuk52zHIFGWCv5r1c5N6K/V9VIAuO3OJSYTxSIHlWy6n5xUUBeLB3khpE
ZzPEiu0p4cHi3CWmfQPKW3gV71mrf+GQlX8o11+yu51RRZ/GqSHCSknvJHzJjrBZCR7C8XIJn6OW
92WRcIIOWrvECP/7pw/XW3akYo2OiNFjA1QEXUiju0eVheAGpqpqCvVZ1KjZzXyVSMk6IFAnZcGb
5leZ1svvh+n/JzW8HfTasEnRoFFJfChHFQw86czYyDLtJwq1o2p683YR5b47jwwP4gtNtSrCBB+E
E3CRBE4jlkJpWBMradmicQRHPH1gDmm+tGq1G46/gg5oqr5hPKx12TjBPDnktQk/REgnFqtmqP3o
cDzeHJ471wm2qqhatYq9Fwafa3fQQkhERTQ+bI4OQi0IoDm2ppyqwK1YqIBacL+hN5MU5XN4VpPa
06kQvvPHXBgqFksrCKdA9pSoMebRiM7VLxA+Cbvl9AEIgw6r24KR6KDYPkfAkxf2+gwHyEbFeQsC
QbgpIopAvfPuTXsy+3Rrck0jrWP0yLZ5xNteQDryMSjSrLDsUGyFo22J8OyqjjGIirniANz4qH/9
PTQL8rNeRJHo6191h514mSv4L+cSOAz10bLHh4H27FbDf7MH8G5vN1QixEyxHyftTSsPWt7sKc+x
ZGBeRJkc8EH8CHwb3RsR4aMGyEAYtm7CnC96hSNm5LgE/2LxegB+ArFNJRV8PqZvntFNfT88WR4A
tketuUtJJFsfxYzjJVBlJf/YYQBh0QwsTn20zG0q8YF0dhxcWUE2pIIs9xwClot8xhT/C+Q+sBZa
u1gghWtMHv1MwddzaW5MqF23cHwX0sJTIBnYy5o4P96g5llggJjOpEkvg8wIbGcak98RSTxPbCjr
JSIU/GC/HsK7YVgN4RTJG9KlSJpsZ1j5facdWbJe6FXhf20C+B3LTxjD45B4YpKQe+qG7+LEFQTt
hvQXFHTxaJWQ3qCtQURqf80oQYBVuIVfG/PukHl4PORHC1T40xJHJ2813oHmet0e3KFrWrOHQp5j
WhRBofWb0sEZ2tWqYzFqTEPQzERScf/huNQt3mmDgPp8qQJo3D7206AwSVdIz1lgKOO8VYfU7D2S
LtT4EjejREvI2SoYmFi3fv/FCEcdScG/jCzon3PIxgqi8n7L0T7WvKFHVLi9AIr2Jga+FZXPdna/
rwIN8ztrMyLaPTiHvzvLFxEv82jrImRCkOAyzemPNnv2Lt6hmONRAqrgcnxXBPXqdVTXm4xbMZct
/TVgM2fr/XDM5Ysflxd74Pg3cFI06cKW3t3mil8jTpm8pxlbzbOso/JEYzpWgZBatEjNMw96AyQi
Ji4MazGIgwtXWyKta9qJa4FuQbIFZRSLDFSvoRIuPKcK5E+RbFiC+VknsvAOE7ivVfhm51Armg5R
/OdlVis3fldmVBPL0d/PRZ3JPatKNqHOO4OaMLwqqot94Wk89P4gAunxKPh/KtJUR4z5YwHfdMfY
GBUj2vBQnka506aSDypW9Ntu+5Z7scfkclu2HLeTO7kV5cGvKruOkNR4ntS1BTSvAsJE7X9dVG7b
dDzErfcyCXr/T7mGQ0N9Lo0f/q8gOvFpli5En4R9pMyU1qTt8CTrtUkZpiPhSkysXW2vpKUXwA+z
sUh8uuPpG4X8wJLzIisTbZVzGWw1E30U2dgOGZBTctcd/kKePfmetlEyqSmY9gapWgPuovGLR9t9
CbBsziBfz0Zs5d4BzJdcRERG29B/aLZd8gcBUq5Ra8yL/6SO6Z2VQFBv4aemBF4dz0RbtAJIJ8OH
T+4v0sF6G9w21fz7Z+BqwV7NNDF97tSQu/MwawcsoStU6PZvNqItOSLluq2jxBJrCkFpYHRhkm2a
6tVzBKAIRqiPjgecApLPxUt6LIhCRq65RX4z4XonY4SoG08vwsUSDSBvKnVzTvRnwRAOsTPFjmJV
EEDByuaeFfyCFbZQYATB2aOeVSSVaAIW9T5Q/LQExdAPTlyti+CgwEb3AqW/4in5Kb7HZP+ElHwY
cQySMJgl5dzIQw6xmzbJbgwoZBPa0bMUD4AJCAIRraazDGZIMqJLLd5kqWjb3bkU20TeNzSFriU6
M84Nt+LQddzhVKcVtDVbY+h/XoNO559a7hfsQ/YuKV/xyz4ISWYx0o9Uv4S+mjorxmUgEjLo0mIK
zriKrt2gZJeYHhUqSNjvCnaIvIObkhUQDbel9ia5zdd5/YREahGBmChth3grmuJKbqrcaWvP/t5Y
dCT1PtdMWQlkj4GqAyzO4VJCRqyh++N1IYxs4jYokVKoI+/sGQ3lRo68/ccVJkzq+t6CiJSeYPKl
tktSayFPT9WrhxOVUQTEjBd8soFIrOZxjz31Zyr2qJ58oLwBUgeipDl/jizmEvW859//0xBLU+WH
pEw2jp2fNsZMidaGb//xnBdP9QV2ESOFikOKUY9TnwXNu3Fw73oXzU/586njyk8M2fH6OGBGmni3
mXxpPQPSimeSVoJ91la+DOsYEbQ3ydiBhb8ALUzzOKrKWmncKaNfVXjjXE8GNHBVuRdjY/HTQK1C
l6bSSvxWTsVhZD2eYsYREGiuU33wkybbfr9qXZuu/Kj5seBzspFHklNsLxs3vA33l64F60uk9BuM
QOj7tX2sE9L3YFn1yEz9zQGMoB97Ies62HEacyq2Wx+pEeYCJTv0lw/fQrVbKbY8JVEi7DoiyMC/
LBjG0cb3cxeohHZW1M4tR06bWfTwPeQVdf9ua2hDFW8vroakFnuy2Q57O5MnHnFM+yXggue35wYK
EnRXYYjjtYgGZeH7TbxGgSt4mm5KRfUeEfw+rpLIc4Vs58FeJDTK5F9A/qndO+IikHBPMqZ74myA
8/mUHfzVu3DAWQcYvFSF82K/x2K4Ohsa6DB5qTuaE/4Wac2fKLZyLloxT3W82kVf+eD6jmh77X2/
1wsGqe5S3OtUk6IS1EPa7cg+avX6dkkCXvHNsi/av8gJ+NbH7SDurg0B0fR5kwYSOhkyUtQv7ohI
z9cWb2e1CZbamlHpfDZl/TJHqG/IW7X8/MBQzwQ1luVNjLiKBDdc0jH4EU6cQegmJto/7S72pjxX
ELa+PL3Z0AQYeUZkw4YzHwUSaD3wuKYIR4WyFCHDjcHjKnnU636g/Lats+m1WBoVNYtke63Nq6Ii
ZhfQYurlQyELqWsp9BKZBdte9Hg/5hFoMOnYh9CWfCUr2S9ZIar+IxC9vVLZnAsLPNlK4wd+jeNL
WImSBx2azz1zUZD/vHgGvm+1TkmvFSXRrt6EJ1PRumUHMaQZtK/pWleZVKl9tCCRcX03cz/vZAzg
n3DmbpXhNIMI1A/vbaBilzInZ6kcqGZbpK0KgKoTBlTy8aYVpEazzvwilHYVQgRN+Sp1p2IYHNkj
Mg/hslgD2Cre6yiJFjqOWqpp72SZ9ZStbnFetpvDaM6MUAHB/rB36zw3mZMqmoqxQITXzAqQdXtT
WcybZKPfFwiBsl4KjoQnsdB20RFx406EpFKnrCntNo+txbJvwaw87ybjsv5hjYG+qd6L1EqC82uI
RN0fFDvk4tz3SRscRNv7y0t6YKutt/c9hmjPsFRfCa2FTElWZ3it/82IXHVZVgG8Iop/Iy1p0gIp
pFaGs+QzU06+wJgw8A4uP7SKzRjNgF2fC6H3hHBly3gaGwsogA4NhB46hBIZTlWknFpY3nNQdQaN
GYUav+hLmwDsxMQKhuItW4KfpP0Csad3rvITFAWr6Id8bCHXdLl4YIahA8bZG6e8rk2QX6dX/LUh
ZN804zkgjNF1NLCTlhjxT+QZOlDiy20a2R/jyIjcTQrGjHuq/GVtPcX2qviPcHzQloi4duz7miGL
qpFVcjOwZEmPXlcxbzGj9jEo6rrxEOVu7aMd7rde6GoxGnWfpBHiSSh2Kej/4GVkJjLIhAK8CwT1
hYW7R0xhifdqLH4uAg8tKiq18V40hMtK0ZD8Ps7gEE+JQT8ghhPNlP4WyDQVeCj+xhxPECDE0816
4wACYJsdoNCMIUTtKy01B/gbL5r7QpbrqjfuqkUMl4pv/d8yy/VxWBpfmapWLFiZ3/PbKPNG1iV6
LytXwUpSuUlE22LVjbumFrTs6Tsli6pYZxk/GUgUY14yc9gn6AhgWPCI88vv33dab58Ph44+MWXa
WgpME5+bw1Y4dwssm8/vEmuV/cT6d0lVdQm74J5LC0pkIn8SV4S+rPMJEQFXD9w5yIXW7sKfSHdk
cNQXkZ2/w+W9D6EnVXOvFiRIrY4Yu1kWXUlcG7NyJmTeqf9zX2hIagunHuDjjWDjKC0WprdHjki6
WxN2kdnojp9sJSHc31WBPRFK463MtU4y8DQQQ2P2U13M2q+1HJd48rHgNEvxZHTh4lVZFLu3Q01z
8HyO9kYbjUv/jZSOIfXjNHp0U5XpP+U8Gfvw3B7Ox+joULd96NFJxCv4vSdHoEK/Y9vCEdO0a0sF
6Oe9w8ETQKGVIAtZ38PSJDlNeowlRzzC/IfICs4FEfHfI65Q/7/JlRvdOtFwgpLlmMQeOsbbjAHn
8Lf2Zrjin9EqsPX6OazRTNrpM8QIXzWjmsE5W6t2oKuvPLKp2oyM/J/0JFVoJuWQZc/TI/Z6Fr17
AQ3/c61Cb2S+/uiZZrqpi3/qsTaaBP5lNvldyHtnbf96PhIyM6Hxlw4JbItL0NRFo/xG57FNHmVH
PNfkmbcMuc1bu5csf25n3t3e00jVaD8IKhTyBjZeXzVc5GMcJ8DH24ez70rKxAGsh0PIR8zQY2gx
pPGjGzjyEmCSZ477VEG9GY7NdymBNl130BlVcv5fJekMOF2BTRWOBkqIIZOVvPeMlDYtKM0geJZI
NB6xihBJFlO+6m2ygaaKkhdB5IitV7Hjt+xJiltp44dIVrc8dCe2UrP7EmKo0UPmVV53Hw7cjjav
l/r1NflH2flxewsTKNliMAXPPLw5/A7/BvEQUpKnJwpYtm6JtHXlmMpO49XW5pJ0WlT+C0nxwyN3
U7qhaiKzYP1p45hsGCZ7yHJoz3WfK/773pQbVV9S78jfRZzh2DGhOFijoutFgqFdaVdaOk+gtir0
WiRjnRiX1hy3rHUXCehKD5HGCrTFdQN35O9MkQL6bnagQYypUqNRUPm6W8Gd26ll0QLxEmpGLiJ1
PiwiVbaPpouHofKtz4U2mpOx0N9hWc8M+0l72MtRSIaOKgnP7WUUSc5dXo2Hcuc3AlZhUtQGt8X/
+oDZrWSSw4cLPU43xDeEPTrd2wDjTJ15Zcb2SW90KaFhA1vgU4KIrI251LZu5cd1DRjRteLBZE/K
vFwbF+0GqK7fLqrvPQ6q3lfpjIkgaHu92pqKOWKKbRuLAMMGGwX6eI+K7qauCKC4hqKxetHYPnky
3loAQpp7IVP0erQ4BDAcytwY1xG2u5kcZ8DNcyo+IV+YfAk/BEYdnH5/XW/wndz3KUporn5cNGP6
SUpJBPhRIDqnrp37tv+qbl+GZ6PD4hByYjewl++FKtsLFfv91Rvwqx8Vm/XgMN047p8uXWt3l6BC
LjLdmJ3OnnGhSnoK2UZoh1dXJiyCjkmd4mtXH6pgTInNBZ1VohISPE7brnra0yBt2sopP7WuwYOw
m7RVoqojIOT/SI2jFmpo20kPFN2/AcCSbjQ5JxcY1PDabU1DNJQxNgSkM0TT1H00H+D/iVVpFp8f
qJcPySaK4AHc2j4iJy3+5r6sy2EHnzFjmW2otWb9wHgk8SlA0sKtVLMfAl1+OTzzul/F3mgWCJXP
ge8q4Lbdfo+ejJtXz3cbRBJUG0gEgo776cy9Rxl8iCMqq3QCKKPKCmJkt1ezwNDJbm5IgS+cbQ7g
TvtsPobD9HhqzbkJnPcybr+yhjhucaDZhoBb6LNBH4UGA57FnbmGp4Xl0RT/RsYUyVkryBnnxlMH
bRRJG05KZ2sawbkpoye+IktSwKe1Qn2Etjw3gXaWG7HcUgWJVOpnGJVOWsBXc+aehzDAJQcCjSH0
WSp8huawBqrCuMjOtoq02AQlJczr7G0yOErXODwWs3XGMuMSZWQSsKixVmgGZEGMq4QrPydUjmRW
F7tofg1XxAk2R18dcvpdTN6KVqyh0++F0O6iaNIGsyyZ71GYaAvRf7IqPviDdjBiSfeML0C9/sp3
QGeRC8My684PxmdfVYR0MuxX4h2Mpz05u1kar/apY1dt+i35q71Ym6HQcnNlDDjfe05xCI6p/of8
gbweZmQ8IxDC/0fUEv1pfgiibM4uTGQc2AUCj6MTHROsBYGeukHnuGH52+TW5oRUEk1MXAZf4vDa
l50sLZjQg2C4hqBNVxssybLgzL3iq1CXtX3tz39TQfFNovQ+11RZg6rZrpFB0rlK7TMrO2tgix2y
EsQhC3NM39wBXvrBdSHeG/PGKE64Il4m/1KjDAeXl3DPo5CBZoQQ/JR7FvpfeHnV63IsbMrg6z4F
/vaJVyLlTY4WnBf4N5LgImHXQKBpd0TcCyLK0tCc826flBf7GO5Gfsj9d015cjQiRZ6EYUJ9IRYL
Gfj9gvpn5VRPRmF1aJEox1lWu4svsi+U3VpJ0mZqjW8mh8qv8B1ehijBvcdl9HNg1hQgh50NPWhw
q3ibzfQVI/q0TShTznBauph6lDoG77FKkaB8BYcv6aMw74xO8e2Q8b9cEn67xamgRprjY3wCflvG
hWdqUT28VAIFKnePrx86NuoF6BydDIW/kN/aDomqMZrBgN+RHYlcjkI/tSBxextTfwO8J3hZiWuN
AEcMytbJjEanqgdJSNffQk64OW842TXV/uMYQBmcDURT4QKdbfo6jTtdqzpVwjNQmWOI+bYlbZhw
xrQejl/pKpKI4JwqN5jfR4M9meEpMt/jh7F0trA9W9aaYHWF2n8EFQkKAHW8EMnkmeHcn46uwjIP
lSCm9zvuG+cljQXm8aDUXYmWpwzSq+PaHoeCx8hr/JJREmWQbQfA0m++sSE8V9BzDptSWeeo1AQh
Wi+eu9zgJTeK8jNzXvilG5aP+iYcl5UjOi12YZv9fHprUiG4MeJb9G29EFp/w/nIhD5B3oqAyr8n
FFI3BnKHaeRK6WElrRLJYDMuzLwgDz1N9xXorD4z0Ok1wmfL4EvSlsq3/UkSbTULBFUUaZ7jpQkX
HCAOIvqqVqI9uS8WCYhLo93k8WxmeSbhHLG5wzVcFKWO24Cpd1zwvoJ+rvoc4aPNrX9ZHkjk7rgv
TM63a47CZWk7DeASIxx/lvRDW6vi/O7EQmAWbIWZyf/RrAAIs+XnHg4t4+tuGCcYUSEZgAeocx62
NWtSf7ik20qYpTFNCoXBwd+rf2xZHitFdr8zwnI/2CXnWbT1FrAuyUhRuhXYplvelOsPQXa7+pZ1
VODHN+LnE1oOGiaJPAtk6B8qH3aguZbwpjfKAo+Q0ruVBsknNAOmbh9lF7GQRlaDZMPKuMXESboe
tSIyaWU2OswuMphFwKYuUAGa5NJKKaP2H57uVrvCwm4SN4W2mCHz70r3bVNNGyVt7b9EEkeZjOfA
n4dxG43lDOkLNtg19hPfUDb969mm13LxntW09iX9yt481/LntmCB1fGdD0hxJ1AdanOjRAdE+NOW
630wbciy83mjFbBy3N3AwSbFcYE2rGKEN8/NUOMaZaITPArkYmepmP+YtXqOA7VmD0w6MyvZQqir
qh3o2r8xtjQaDeRYRqYenVvLBaEIrS+xB6SAifW8aKfKFTJDV5knzaMGzWoRcCnM++RXkz7H8HOC
Zq794kJ2mBWMDaBDZxu1+hQYExWHFrDEGBKi82sW89IgHyy++m0lvpzhWCPBASsJnRXrR6aYwldR
RU1nWfuOuCqeCL8wC+RJfDuh89y1Tlg4Rfeb3HC2sQu6UVZKm9MMGzqs7eQsbDQxyUAPtpoFFNN+
3b9iL6NVeZc5gQvHVUFwQ8le6FxrKfoCt9TfyNqZIsRxxRr0pxWDqCm6NHhxeObJPDvpG3C1HLo7
2gUN3469bYY51Y/E21WFh0NYQMYzmHgN3F4qOHM6lUdjkjwZC3V+cWZfnJsiw/0+t6Qr5DEDUjGo
4cLBhcyjogCvxnrJEoPvsFCZ7WRzfBkztCAlse0DOI2Sfz64EI1bleI0LbJGzF6fmEstzPVAGwy5
PnOMg+0o7dEpHwefs6b1grNvNVLCOvZ4m0qisSYgp11w2s7N/3lP93CIbK5jm5a5dY06AE0/7LnK
qGVdYQVwTuHeYiEmloev3mUBc7m2gkxG+KBrJ5epoqiUjJOtTI+in4EnJAjT46s6KlkBYDTQueYn
f5pnXvlSEZA0MNwmCEGkgk/0++wMwq+1ucSkdteKVidbNjuruhXVWcW5l29p6T2yrYP5Tboc33Qc
G74yt3rwNcBJuMLleUuV1yU5ChNdGWa0gZ948fStg6RYJ79tL44OBv5sD+VDdOFWJoBzlH8X4hFF
XQ00pbav57MywK2H2SXdPmPHw4mWZRYvhOxFkEC8b4aPIcWOFAkL4K6RrwNFNl5PAquxdRHWCZRs
1QHp3eBLaDu98AsJ4RN12t2dC4cQDQYaV97lrhUt5Hk6NvoaXuLs7C8U4AzMJn8+MJNq46Qnmn/V
vUlqIOm1aeMFId1WIpDzEqtTxHzayLLieho9phAHiZoRdy7HybKuRFoG8YfF6B0T9pGfmHBD7lqD
Ni9HqeaFk7SHAgZ7GNhvXnxyQFmcUollUnOsWKaNxASpFOj1iez1rEdK8EhRTcDgMtAf32mY1wOl
x9DHy8ntn18EyKgRhnbiuRm18G38SUClG5Y9uibZ4Z7mQMbP7YgYwpZ1lBz0fSPKKvjD7lq6gbyA
wzegWGUSdc2l683n0g2mZjIseY9ELoNiM7UW3cVlItMd9l4XL4iM57pxmkfGJZ1HHKg1kcU3xacG
bJQIz99FVGJyEuLeBqvDGMhq1IkkT+1U43fxDLsG89PAYjTkNiqdUI9XahYYWxyMOBULkvJkcfpa
aFdIes4i6wEaU/esTNRiFPHjPhglLdlBGCQCAI6vvb1nbf6jLjhSoSrpZWnM7jApTqSWU3i9gXzR
E0THADipOajSPipz1xkG8QCyKNFGjgu1Ax5DvrJJnGqjL1njY7dpqGUQJHMfbCAkj0WPrrmiRxOc
HFFJXRElMd55hgif3DiXmS8d5hJPlaCHv3OGXWD0dKCxN3/dOry5tv0etwVs/nBx5flKOCtKBtwF
AS5MaPs58FqIQLMMgWCz4NLyXwRQeCUdqOLh0HyqLjLi2e6lSIGD0rEZCNtDRqJHtZ7c2pkMMg7Q
1jZJZ8/FsxiFjeMFdSpXQi87Rt16UmmUiN0um3t3AdpRkI5zUuHE19WBryahCGGrrtI8Dz2LM937
EpXLLCw9c8bIhH4ixLAdYbcLujLlyPRAGMHqGwqrOGPv8Fx0xQ1uzROzN/2aZIWsjq82ugenpl2P
KYtW9qC+k2sNH+N49yqbifHfYzoX/Uuf/pDsh3SVjonJWTxnSvgt3HgB9ut+mMAF4ujO4rGuazyQ
/4upKmjlWLZq3Qw+LhGr5gSqXGII/S6SCgMhyJJ4Mz3mQTlm+9PyV7kYRPEuncEyoAwt5H/1Ap8T
N76HEDyA/BxQSGvKaFFkK472BxgtGqXtMH1tfbaVfcqNETJwe4PEQkSd9xgm58X+UOTcaCaDzHc9
Ez0Ho3JX/20YCZQrWPeEK+XnNW685y7tc0v9bYNqZ2j1zcPDQgAvLUp2QuYaKmEZzvdXscyQcFGK
XhOcyu0mHm+iTU34R5MJCiG+NM01ZrW3dvlpozFCUtts1LbSWlZpq0KutRLStKONrwGWz4aIXoEV
OkXSev56HIpqQimkJLS9a4ptBXItbvvaWcWJ/LO/hDx/vC/DUoTXIoEEot1UaNp7ubdfAHF8mN7G
tPVlvd8XgW58x02qP8KKCzq0SfE3Na9seKr6muKWBPVU/NgzGSjQzUYypUPkuOfel7e/iWxHSoyi
FKhpoIg7hwWExkyGHuK1iYcSvCltYWHYSpQ20Ki9CSRUrSuS3JQ3vSjDzPj+R5YBxGy83Xsghq63
2ErX9AfSfOXvMAUvXyMAtZZ2rT64jV080zrKRVziVE0aXKE+HzHb+TQ7J/15Nbtu+478X/aa1sN/
cTdBlqW+8sKuHiTYxTgARBbviYPR0Dd8UnP14pYr4Dfk3fa5aU8IzyGAfMnCLJxXc2wPcFv9mEZX
yAvTcIQ8G50kTudRJkeUFTfo2ftwEqPOOv9OjjvuZFglnBTER8iGpEDYaFIZfKh6gQ9BD4o8D4qe
zFBgB3bmx6gi60XLYmVMbiksfP+NcA9NwOkWh93t9/dzk1lmv1PNWVd4VDM98ouf/3w8fiULjW4Z
on0kACRJsnhlDE0to/VJHmm7jHBvHimecJqs/HBTvLTeryD3rxW/mSYlPQIGKn/fRN8IPmXc5nJj
jMSviD3h3tjWBY/4t2mkCnil+k9YNJ1zU3QpLh8yQG9HYycqNQU1W2ZsbkwpFrTS6OAqmh1FUarP
AiOyO5ZHmfheEX+yzh2lTRbUSDiaqIyi7KwLkcJ4Ny/AYEz6NxvuREJzUXlw/9tWmdRvY2E8DIDM
kVbW0xwfR+J0COKg6IMr5nYdBN+WNQf8XErEt3E36qo/HCbBZc6wCblM9gXQHat+SK74eOktEv1K
b0wXSPNz48aJYfbUheU0c/F0ffJRbz2znrDYnQvljZQAAn5n+LstwlwLXzvfUNnx9xUOz5cMYIhb
YyZs3DDw4GKPVUkwaG8HtnxC2VFNu404YaugYlptdyN9bRh6R5D3VMEV+Tpy30zEj35C5C75mXh6
VnBie9KgAQJKsmVhaRKEyqdh6x9lq1so2tB1zLxmrn8DYRt+sq/IggilzASnjj0JS9jyKhWkx0g1
BTG0zJM2FqSSXRl2SiOT9Q2iggVNV3YfKAFEE1juTZXdOXv5PtNNPKDR1AQ70aOlVG13e9ln0QzJ
jTRyKOlAfNDXmy3ILoN3bDI/hc0+c3jcBXxSf7nkmp52Cx3XsHkyLQqBeUkS5YBpdvhuQhID2uXi
Jx4areULMZbvIdRRN5QEa3UlDiLi+bbaNehHWvt3G7itp5AG+OL3aplP/64Ak3/2QvRhsuKW3AMx
+v3Yd4Gugofd7eTYK6S+6sTXwNM8vQh4182b7cO2AAr9R84Zt1Ih/auQWUzO3vD/bT8Sq2BE3rrX
NexmdSuEdHquwWOrJfC6hORK2C/b9nGMLhfS2ikAxCM7nW68E8/sAex9OVrX69gXryL5JMA5mp9K
Q20UfRJBbbx1fzLnBBb6SghCFvGfs121Tm6X11clcILgLWGzrhVFn89vNZW1YRLKLnUKMByZdKk6
igE5SqseNN/FuRmbfDIyqoDlcNE2mLMQTp44eG/JlpNghWVARFdcpMdAoGzz6zzzpARNFcSFTazL
tWXSJ6by5I3qC//ObqlV9ectIeMgMJ30WerAWooeXfFfSWSIA9ylIoDMrtNclB3eMVWXb7+ekpql
n72rUOCDYFwTxGuKKyniIkV3Qm24rgkZ6NZyMf2+jcuDNszmuixjwYirS+okZD07O0zAnnWp7xsR
zqm6OKEpeCdXgrUqka/t9NXOe+fpNXElmVJVp7LSNe/+N883R6S1Wgg8lTLGV1Zns3aV9ZxMjK1b
2jo/JG6xnmFpN2h+AOJ15+81MbAlGBRQb9RtBD606WKsjPC92b5++4yF/HUN75UFUG27R+4wfUY/
q/JDqyD+ZN2+WbKnFz7+teYVW+zF+mUtA+DZeD5QTIaVjZNGcu6EWazE+KfQdVwHG9fuSmuKTAiI
5IDVvTHOVezj5/v/wvbDGcHAEwXscQkZjj0KDicvCOOcphglgkJDugQiZq5V0V8B+pcTBuUePqK/
Bf1TwWYWzYohU1o1541wrJKfaZxUCJopQIpOzf/eWbWAnnU2RvVM41c+ACIQ34VMxUeuex9O5fCb
A7ZxYwqK0Kol5FWfApb2OS2el1kRIwU3u+5N3ERySDWYH4MyZ8J8cvUaHlH1eOo/YK3e7pHN0Md7
BOKrTo0manbTYnCoeUZvsT1E+7DfpSCcgqGO/qqotwpUfLllFalP6Vf/8N4k0AgL/UPfz7mwBQmn
txFAR2RaZqeztlvqWwbvsuFEwgMbmjb1PgddfOsChOhB9FFXQ3Uec8W/JZoqFikFNOg5hSWqGFba
bdaVR7bbCdqEslD2CCH0PS+fVOYHQFI81MNjTkw7VBUHrY+Zv17cN2puZqqdI63O1PbzCbCwoK6F
CbcuvDtkMoi6rI7kibpyXS4+AGkHhOgPehSA7V6izjzY2hJihBnl2CXkPRjzwlcguCmvTEAUqUw8
epynRdq+ctiq9b54+QIucy6QKs3RxRFzxAHPpDCcwnhCXLRPHcY/CJAl/f/du6YKU1XhaP+5Id30
8FJsi8ov4bnpSRhivg8laWWNhiG4nMXos4XSNgtdvt5FCqlhlyOOrUad2q1AZsGsoFJ+IcMzsvpH
csMj+MBrjynVvJf55r3uVpBLsBgEy2UXCZyKL/XYWIjjbkI1K87W65GS5r9erEPaRV1S6rcmdRz0
b+ZXpspIKjAKs+WF+U6/vBaRRxmlK9cbXUDnqS9vmnVrbncPM/lNCuEcVAKFb+pMqO/0T1fMT2oQ
8ZgdZp2kjWouFO/akX4sojyCpWSzlL6QY/1PHYFSYnwY55a+AiLMiUPtdVzqXUFO8p6sODlxyBTO
SDtMOyZYon/oIfqXNCBoWoLVUvFI5MFX0pLeC2RJJkZ14N4Bng91infxApL05mduq9E0WK4M8fQs
F1bgSTCV9i32uNFC4+/SMz4cVFn7lgHF91N8Lr1D21SmKH6IVWBDM0rX5f3+05NVFwC5vc18bq5L
w7sUNpyfBhyPmwE/z3tHDzq1PoSitqCI+PAQFRh40Dy2+zt2xtLpql76U4e5gX5xMgHLUp83QFT9
2mYRAP5Qcr3JgA7gQApNwZ8/48imRJRYwXcHXirSi6TPLNQ5UgnXj3Uu8KzKVlR3ROOjTmrfo2uQ
rD67Hl6ecPS7go3g/BcNwNayjpLq2rW5yyhG0dubDO+abeSwf26mUhPG36a9bzc2SufyYF0Sw1WH
1Ng1NsIsZD9+tA7jH05DiixVqUOkteFXMZyPanlNOyilEdvfglGQwbCSpRTalrlrZFSQeh2ydE0X
Mzxjn4E5a7chKUhaN6ZzCMICPv1PYzMmF+LgZy7DXMuZCU7DawsToxLbIafpqV3UB106d5FZPyyS
CiB1aSTAMhpq06ZK9H5L50QKcq7iiTnEhAhcW67zGp5WlcsQgO6Lrdeiwbe6iOlHn+AOKT9TqisD
/X8bVkddFT6IB8jqEwIXLt27Mjb9SU4bxo+r3A6/DW57jbooF+BjTCHk+sE0J2siLui6rUtqOLrG
ZF0dRzH9AQpNRtSPV+iCcxTQDWUko6roMy+LRkx97yOAVW/3Ova2QSNFYXRpPiUVYO4+DC1z5GNJ
Vfi0tmRmYBiOnBp9JX6R01hGj/2eSmwogynpmSVi2MKDYcryF2gSlp9Jzcx0dmSFxoBxQl4ksYBA
tn4V2FUUJ1BhharKSD7CqbCyhFqkXhqbZ6dd3OdGzDbtWg1EqYyoItIRKlcqVvU9unvIkTwgaN0O
tAEAlkTYRFMTNK3OgYKu3DDqTtYXrLU+B0of4LgCqE0+Ji9zLLlWo0dGLNsUyZQibAD2B914e+Xt
tZgNJwbVBGAKW9ivV+chFHkPD9yueb0zmv3JswloI9Kb3C1b5tP2+pEJhqGmc2egXMHEG4dqGw3S
c2j4SxwOLlMl50Xe2sQtX/03Lspl1sTJloKCEDcKzoUT3pmcKXQ8bf6SKhD2/sbTDiZx1y2K5feg
kQugO1F00QzhviMh2YGaBf5HbwC6dDEA/cmHbGOhaY7HIsy+ARlx1TVnBAIWI8AuVycW8e+AA/Fz
76Am+/rxlmeMQ1g55NGH9EYYgQsz8yNmCMMTT2jDMx0BXd+2V1aEfdDoTh1csk+0vraWSwyLqyZE
UKWeTjEczp4JTr6mm+QArP1xfgRm6f7lx2whVDOpEdrdGF5mmk+NioCX0JdxvJxH6w2+yjLcdTRE
Tqxp1BATmH5F2ZG1KPTskOKfCp7rALBWbOXhRK6xGakOkXpo+zzBYYKrfvoFnmKEqiUMRyivRD6M
cKSL0cC+Qc0YbJYWXR0V07Y6sV9qjYtw+mpUp5Kn8P1ZRHn8kU+5OmAXQKy+YqdYTHDV3kdb9OFa
MKpFhXeOPOXv5EkePUME212/YWDv2qKLY4fRFj77It7D2JgBOaZmZesRqumGhAABpbiV7J6pK8qH
591PxNIrLBy16SCqxNh4+JYutDkRf4yFUcYETIzMtvLaceScs/wwLvtcg3dmHwVMnI2AOv0AqNN2
fwIkZ69IqkKGcvIHfukfJnO3gQpGu7FGq9VvrrQGWFKdlvs0w7y3086p+xVznjldf99WzB3m/0KR
7jCFTXwFvOZPYgXurp9SUaUx3Y8XWHPv1rHg2QjG1hb+4QbxflPARaPBinEvoLMYXORd8IW3Gf80
gPrZOotL6SupOnmMchl21QEb5uJ4E4D7T7MHmbfZfDVRG32JqrK4L9/QYYZ/bfvsptYKD4u6/fEh
4jzPKMDDqbMHFKD4JuSCpaIppkJ6Rj6ySSQ7XsJd+zgIuFcLk5s2TJL+1OqD6n1GA0b5GTJ2EiWC
NB1v3cIpNQu4Tlw5QRlbu8bpMjUUuy1mv5/VWSKdtRhZ3MsZyvUMzDJHDUB24jqJ0le+DUbL9RU6
WzQwac0kC+a6Nlvg8z3ur1JozFvDxOJsTQHVt1O6GG8thD8sIs2F1+dWuJT4VspKJAcF6lAvMqZ7
D0pFUCUqtvrR2qYCRU7HnEnBvsJDtBlAB7gQ76dbHl3KJNt1Pj3ejE0uPMY9Kyab05+BqarBprMM
lXaY/jQ7nRRlxVENnXyA0PQt16yGo57jJ+BhSj6IP/mDV5cXL2D0PTCxDOKJTJEBrIk+0aD2pMEX
m3Urm/aBsDXwgPlIeu8ivZ1p51dFj/4PYopDwPXs8TdvzbT2v8HB7JEtnCFMjNgeeoM9tpfg1V1l
sTr9QpwzTcd5YRpSh1Alu5hus51Fa3fjaz9Xlc4pfRSLcn9XH0JOBPLv0ohmzcAXaGxy5DsQymeS
BzI/dlvJEKGfwiR7fyJ1a6AUTuoxtt6Vu8NGyNOM8A3kHtSGyPUnSDfBmXBx69kDZUodh8EySnnl
n2gtQqCNhETW681xNzs5f6qvmgM0oAsgq6nqJw1qC6yedfaYKngTbRq1goKrgrjAk+dz6DELasDc
mD4ou4PG8t7eftmDRz6/MTFTv9XsSPL4Fr+u44CYAtS8CN9KjbCxrsMCb7djHfJyWdXgOF2BaEWr
VAT+R3a7tdX4L380NT0Vlk8ftXySsHqPA1Qu7pqzdLCLt74KFK2lOfEskAgejf8feY78kEjGICke
w/N9IbZDc+mLblhDEG4CDKy6xJ99rFYvy48GKqjcmj3+dsvDt8h8FnpCvyNENVAUWgSaL2/Y34dS
ZOzWakNxYwqvd/zB9Ox86a6crRT5fjHqni2ljtpNG+ni5pP/Dz3QyMoGGsC130f2lQF7g9gNBEkG
UNkRJ22KYbK0aNIJ5sEGVfbAJP6KLJzP3+4kuhzmIporTx/YZRZolyAyL/xRUCFVjs3qfxky25Ex
yvwQ/KkElwXAWH5CRpq/t7d1lcHkLRFnFxX9mC3HSgQmJBtPmIyZsMwq98bMDK1BBcnGWay17gLL
7l65RUr5m9BXYokcY2Zc1/rk7wpKqiBvAr2lTrG8igwK7svDYU8erc8qo9SiFNvW8hLpJ8RNO+hO
pwU4zBR1ZvqH+rd4QdZkvRa7GQ5iJiI2BY9+pagzsa1qH45RiXMbX9VbxeKu5KTZ7KW2q6qZRcni
dMjontLcLrD5uwo99UOlQ2MztLG+P1inYXJZd5d13UY60JgP7uqEI/pRzHq42GQqC6BFc6dLc2kM
5u28zE7DDFg/FUil29yap8yhhd/aQdSswc4uOnLOXUc+jsWEPlf+r7VAVlU8SKEa/AkqvT52+Dpg
OwlABY7uOYfIyl7XhViewYP8bTz5p9j+hs0H06lEwATFudz94DA0FnLnem6IWqVoZFY/97bl+vq+
/ROuhvd9/bQn4FdHbS3OsSo/VyL6BoqJNAY3rUPWlCW0KSUDhJz/9TMb6JUE5POa2y4QpAH1ECkA
4j62E2yTjkd+ohYYef64JfD/RUJfFdk8RWyly4AEp099ts8AS7eiiIED+T5HcZXXB3iRadbqKwKy
8PwPaR9Km7wQWedcli1Y0mUz4yj6pBANY3ce3OUJeB/tOtAMFD0QMYI9CPjJrOPfc2BZawZptFFd
sreqUBKFXB6HpD7cgl7xK0CLIeFjb4jA6/w2BMNfq/J7NPbXAPdMjcjvjEG4QHDBYlybHvFA97nT
q3aMhTFRpX4yyJRbtTX1jiOj5sUj3SSpZ1giJC0jl3LUNFqODvE+ZnVrcaAT3HTjhrgbfM73wUAo
7KE6H8Q/JS9Iz3IqhN9n7WhFjig/Gw7+bAaaK54xsAfMrooeHUXDKSySNq76rplHAGb4cHc90WKJ
cADFWLi61uITLe9znEISHp2XTQJjIevTuIyWJCW9PyiXzbxUcagJoAjq08HwRIKyQs5IxlPItQop
8gDjNaf+jXjom1aA4PHbAwpTyXV2VD5s9RTLAM0iM0QH8FCxF8+g2UczblaqBK/GR7DwtL4hyNIe
yosunSdeKHEHytedeAKKS/QC05w9gz9XXkpxU73Ws9NB8MER9f1YO6ggKTeZvb9yftrCob9eOmHs
3LX38IO6zWQ0kIjJQANKhSm86Sb2l/hSlenxMkrFsxEn7LkYnZkd6GVGo0dfP/WflEKwxoVTXgT4
Zgj8o7sY8dCDy2tw90l57BKlVTmPgZX5ddHdLHmQgDlAaDCXm5t/xRL9+syIZQMWt/RDAeD4iteh
wU/wi2TJQbmXpcfuHpR3LZ+sxPwMbSMQwTdNvg2YQagbFKFUODt47lcyAewJrev553FIZs+YZ/yf
A7WgtS/arkb2Xg4WIG2onibPW+R/cz2xoHLoiLH8rzcW1vu3aulYFqdHnaOONSizL/p9pAub/bOh
bWJicf5VONcSW7ErkJfp2UqH7PRKH4/DUzzxSPdFCqHo9vxxTxU6J+xaKu8zBWiKnwiU1UDYSAQG
0ESAtX4v01MUBMSyOCSCVkKK31JhC6Xtn7YEDcFoSKoqXcwdf/eaIznsQ/4TcA/Cpy+FnDFDt+tN
AecitRs++Alhs9G4GW7ItVGFhzf4P5a02GTHULxQhfWYbYzyhSdf2e9u43IYqhob6YEhPwjoeS+p
Hd7OH/CYsXAVSE5Qt8YdfzDhXDZ1TBhA4yHd4BTaWWbzntjt/qkfTklW/Jb8zPCCv6eyX4bpHcQj
04JhXsdDGOCa+Hx6XRxIsz8OMvgwOwD+3jjMm1T2cB5PmfIN9IxlHhqyuWN4qMN9YveKGegroW1I
pIKnSbEurRrYxemXdANOkXkwXFWfFNkYMMY0mM7K7rSZr6c0M7u/TJyGvQCz7dDV87Hj7KnBD2JJ
jVjJYG8BEnUJbUw1Sd/ix6gHqUZfHr3gOuyhEX6aWLuOAdYtq6Il6dhSrFRDhouYMKAZ9/TymJr2
vTBDJTpsTQxzWbxMLOE7IOrVgx4LqTC+nOLuQ5rJUBLMsGnYwD/wSO7nqVcisHvb7ksaNCdmHOnl
tYt9GrFUXLFwA8KQ0pvufoy6qGmP8p4i1QT9S0IrjL2oD/d38L75ZFyK9uYvB1TA3AVM7zYFwYh0
Frph+h4aSpjuUGXOQldDIrVOmCiU9XO9aA/1d+CdfIQFRkkKTsEg/GaJJMc058Td6X5JwD9xicwp
bEJFTygB6ZwaIewA7zNJsj+uBeiPAMkIlYPwTf1VsRjrRqDJYzznxdR5EjUmMDwyyaTXphIiHpZT
Wb/cvnFfiAIjv6+xW8opzUjJ+7eNiVCm5PTcyy6KfmmBSnoKsl741yyP2OujNn0CfXNZt9BbpYa4
VmuC392mBLQnFkPcG0a0zK6eSwYgnPUabuOCCK6a8QJynDKZODUkomAS9yavzwOglMtam6npwCiE
fCyhhc4Drsg6VZ0svYeYnmzOSsqc5JxN4pQOgsZNQEcH6TpVBucR1+k/hnXzLKF62twN5dmM3rIk
/2Qvh37p11/e/cKRkIjOs3WBGKxf3IuOp0LnV4BW4nDXTlCRTO4sFcXVqjodyeVGAb2Xt0Uz+4n7
HlBws+1Xo/Gx7d2MChKRb9E8vDjRYFFi75XVH+fU/NAo+YR1iSiloZli+zTkVMdhytY8uPeiTGHU
9XpIB4tACxRih5UbguGmICZosgeciWG2VCHq7jDfDKexoUmIcO3IV9GhpItYO+vLlWoLuxAwOv21
SiKHBY4s8CGGycsrq38Z9PEtj0hhARNscEVFvnmM3UAFkcxRY9LP8AFHaN5ofU23vvZi+xXcVIqO
wZ6br3nDQScDdwsYgNWAnIGVD4G3xWg+hHkx1qMAdn9qxckLYdGjzJ7qtjCsGutPVd+TrpGN810y
VNh77IkXD8fDiGijFQxA+BEv2l+Vt3N7ZZsKiOPvh+FJGQNBHqD1qCpxXbD+U4xsecu3HDPnpM8I
zz0by6XDPS3ncL/hIuwXhP2ULo6MEx9qD5hVHcsFlp7G6YAFX+9SJaESZfAcMD1a88rcqg5HEMbL
Uf1zdcCwIAcavBaFBCNFe3eDwN57ofFXmF8RBAKCPZS8R5uJKh0SmasqL1L/VppntQ+5BcsqdavW
zy88GFj2ak/PCHNjFK/CXJEwDr7fryRMOls287/mlCIFdo+QVF6yOOxFHadvK4OK6NvxWKBne6e0
GsRTJSktTx4gUbpf+kr79Z1iYXUeWbkccycXuFes+9VwnzmK5jO3IR73OqiAAaOI8rlVJprwEAE5
hgk44XmQ2Yu6fXKZ747+lnxUnX/Gupw3Xmyx2V1Qj72FxcXJU2/3AkeTHK3Wx2/va59czsGqGUNt
beS4zanQEqtDLFIDMZyIkRWrJq5oNtKLI5IBhmGqZjE/XGWDTiQyQTvFSYM5b5HUuiGcx6sdOGQn
QcOqeT6Dk5+qW4A55oBRAWAod28eLE0kx4dRn4Ye3Vgp9B6HKRIRbQUeQpjlHy+Tut4Ih2x42G6P
XNkgfFC4qbOSkmZz/NnBxr1w4AhCPJNj0rclN+sYAW5Qx9oTy3Dnsj4P3ya6TLGQpp4cTVVMkQhG
3mLFYIi+FMVfWiOMVzEosTAIWtXzKdi7JJPdeCaLGYG2MnsKAJ8UMxlXvb/YRzjQbNr0tZCR7F8B
Kfyis1mQwNuymY5bMJurdxqQfynNbSS2r4xnPbJCiX9cpQxNiQUT1mAZZVwoh3GPsJGs992BA6GC
OdZ1+8qDF4oe/8wPWsBgfiMu5ARJuszEjgJlmjJvMg5vJQmsu3z+m3g9Hncu8dd0YgzGn3CVbEiJ
gtxsNSG/VA0zl1n1exsvBoj4A4IzxPMy1PRwNA+2SYLmZljxmIvyS8Z5m11pCxiFkqy7CH5nHhKl
ZmYA6Oj9/oMtWG2JceJePQAonBdXe69Ay7BgUHWiU8ekL9eEU2mS+EN/1iXCrEzUcJM2rxrfYC5n
eWTwyye5bHVj6IzTTF4kQECcerPMaqq04ZHbceffX3Vl3e6y0G62CHHKIzDonU8U7tpxAYl0Izsc
jv5IF+ao3SQadzR/NhKpnqKM7MfCw8kYDG5yTVStD3DxRO873yRWzzwKSeHR34yVcCjY8du4H1p0
wjA46+M1owswNXb6MAy81M8tS7w14KZnwXGOlhuy/Ikw+1k/XxM9kTbe7VTAJGGs0NJkMch7+fxt
9yKgSAURJueRo/kmbYRfI5XicDqA9OOIS5Nab9xNdrGS3hvVn9P/pj6dxG8iOt1yDOaeUCaLA0UI
kEcmB9JqIoJTgyzV+EKggvMp4Q7KfYMoH8omzxqzC7Lks9lahpo/Gz3+VqW+M5p3PO6QFsDov6G/
8o6hr5Fk0CVuM8uxECSbL9CIsLnUyf5NuLhUbC8u5QEgB2a2m2IgB6Z4iAjoS4JZOZPCQBSm5HT3
5iY1UpP0rUfINrsV7WsrYbOtiFeyrZydibPWavax+MVyvN+bWn3UrNLqynXMkHlEl6jaK8vVWD56
swuPzwGIrMv2y8Xr6bjpNQq2t5KnDsmGBX7PDZotGjdKbtByU/rUVJj9/CAUJBhRminReTTTJ+dK
39GmA9k2GyhvaJOHJ3O+4LHBwWD2QyB57EYICUL8grO7Xj1qJuuNnLbgaENY8zIsOgubt3a8Zd4b
N6Dp59G+3j7o0Bs7ij2Tmv2ZYfKN+9mkXlUsvpr0t0AvEiPjfSzKXYzgj8TEhFiPQXrXLLbIbfjw
LP7MBOhkU2cc35A9HaJdaeZeUXpuK+ufK9ci4V1GNTqBqy++QsXvyyyIUwQ0PbZ/hvf+Gn0fDvda
AXJWWnaLItPaE1lZCnPyq3yeCvtZ6s3/mGQ8C2o8VYIYZEYBnxMoKkAu52GPKjOUSZ+APxHCtIeF
HIGa6IJESVMiLPP+4KpYmZL9gzMeIfBc8cWlCNbRqxFXMcRQMU+9ohuvK8CKvpcl4t+uiit7kPBx
CXbf5upi82czxh3RXDseZUAPqJfK4Hqeptu0mckfzmS1QJRLizZE4qv8yI696rBR2gmhyDoDrval
tQx8F5B3Sb9TzVZFUMMPnjXhdmYrRziF7iQddQMsVzCbdki5HPecXUIZem65zGEddEDsxRPeNGnh
FkWpTrpRuTBdCK03y7nZpTVvzVZ1OLyDz7EmRbWmiT4WyNyDArZkfcPPzhNYGgSLobyVWa++P3ew
JYcf4kbhdFt4OllYw5vhp6CnQjzcswIF0MN+CsOYQHz+7dfxqvBXOb8vRKTFnQeSmcMi0o8P5mcY
WHvnNP5AhAajpA3YMgB8ioXQiqb2CJTJxrpjCL2AZG9oiBtSIQNP4B4QBbb7v1uruV/ykm5HO+O5
6bu6lPV7i1AlgkvqV667tRPl37ccfbjKeGUukAtfjK6ORSfJ+BfT/CIJpTSUXene/C7dwXXgO8y6
FHMoxi0Whe7jXuNyjJX1+hfX1rI3xjmmhLadwZMwS4vi30gILfKi7ymmKaOUW3s3bj6OcMjLcbGy
+D2oVAqkCm1uzIt0jt5QzYuGRjt7UUO35klkGUpeBiy8H0DzHrjiJFa5pfATI4YCJsV+8IVh7Qi5
QoqSfmO8hwHC9N8fREHtJmc3E3BM3F9jouJxQywe1WwGcjxyCSF2Z2y6kYmqlWEpCQfmJOS7u7kM
v+wT3h1j5eBQSW75ruyNizcCQjntux2xjT0Ml6PiYaW0dkjG4LvukMxslN1+Mdchpgvui+ZuiMwt
+5+7buXf7HC6pBse5rdQtIkcU8gI+UeObauG/z4O4ABuPJyIQ0xdCmUO4Vy0mlHU6k+lpeVTf043
pRM9HwhLfPsDJ63P//ph0eaGaQfZUHWNQCX6kKysdHnKU9+43rabgOY2UJpYR3zjtLB6BMF1htu4
0e8DKGTR/VX5D1x+GVU6cGhiR/iIUts5H6SF12rBEf6XQmvzwoUQ9s1cbOJMGwBOJZRaVW5PVOCX
nnrQ3PH7Op7na6wtcuAovYzjiaVN4RAYz3cPszqs4e0X3EJrzQhwFxZphxroO+3dzF9UrQ0et8Dy
zra3MPJu1S2bXqHNXxIZfKOUTJDjA2VphoFdrsM9WZZWFIs+oiE6H6NDLJ3GwHcb8B3OLlYx1cmc
xpV3/kuiFNQSRN1/xoqI5tzx3xwfH1GinAkIF+FfnijgUlXTvFwYvuHeCr3qj5bRUeNRPHY386nF
hCoUOaoz4NhLSVkuuTSXGkZXQl9p1Us9LQsucOGXkEyB415X9rNavSRKJN6pnapiCYEYHE6CVrRv
JRZaadm+zwTFkKlhs+ttU1jlNFHHm2OkswfG0yp1/7qJNp/0JfWGC3GvYWuNiJ3G3j9ijmHHIROK
Peoby/ux92exRuvla2NKJySuH/1Jz/9J+2kWsRKXVtBjtgn8Wh0XXwADHlQNm8cnE8kYwe4MPiu0
IjgKou/05QnKFGlHncFkdUqWwpeo+LY/dYLUSj1hOIer2E8aqNvqAXS25swOWgL/eIiBixMDA4oK
Oi811p9rN/ZgxXh3V4weNB9lU5vSj/ptJL6KsHpWzIRXnPew8DO7ymlU3/aQVZQBPAj8xixIqcOj
JK8qohpEEe/3Tb0UJp5QXW8OB/g3g8exOrrx+ZzUs0hMlGKd5/RTI1jPTONJInazhtcgvOfuXfth
EQDtyH98WfyFVaXRwq7ktFwALkLKsdWTLyUabLUPFEcUDghcm8O+jx+FWEkKToTJntS1PshCOAgT
giRLh4fMJkqb7cpd/aQ7tj1+8xl8fkcEGh+j1XrwXFppGWo9KwQMTUZUv6RdzKJNJiN8fTeEyiOD
GPvanwEcWOj8kJAmWhkqlTuIeylGP82G8FRfSsv5ELuFSke3sptuZkdiNfzi/KvKHpfV/6JcmDCb
+2mePP437VUBD07k2UVNPevAFCjwIPSOe9fbbjTsKka4sEZICtO0kwaPGitCiceSE8TjYmahYv9e
TSZ9kQIojQ0zShw6MVpPaCxm/NSU9QmJV7aktEE+lei79OaGMynq+NC6KLfn+Bk/idGa5rf6Ojbk
1CnplGk19hfQ6bOALAcyHd7/LYP3rqdx+VyIEyGYadwVfyx3SZhgBoXPzwOBA+bQAKwNy9ZjxnFZ
meS0nfLyvvyAGkhAWHFHmpsaN3BFXM6BUaN9NuAbuuT+yLREd6KqsvJUbnR/msLh3IOsRvfcEUGF
2M1T5/VEAXo404rEuf9UYXou1U5Klty2jm06GmWLyqAgeTo+g+U3A+KpgYtB5OUTbtDn27obojXE
6j5Jfl4Ftm7tDh5vl0dfY/u3KlpFDm1+VvLSlksaPomc1XnC2zc2MBJF8fRpsedUwPky5yVJTiZw
0g/laC8U45mjHeEswWWGhlgMRx+ipKHFCi8c56pbdXK1Q+L0vt0gHWWWUPSxct4tLHoqCzP4Oxqx
Bq9mR1+EW4ypyAovcaCoKmRZ/w3t3quxaz8bjvBFtvYJfxGkBGkLH2fw0hgRxVoVSwLj6CL47HXh
cM2lIHHZhfFBoy6v7iM6+Q0tW0qAPgGxbknuQJGjoyGMU6Lnm6LFhvFWmS04a9QJlCIVOpHAjUIB
B6Rf73Ot73V/Ae5AuG+bAClkFo5YWlNPq/4pLZJcvxoj8AynVwv9G1zAoFU6+W2x13u+YJYXd8UA
U/WtBYrVZRRaTesNBqFHhhojvf8UhOdPkWP7y6dQdJP43WLFLS5hqDiKHHJjMTk48sPq6du2JzNc
cvYG5mxoJlKLCnDO/AR6cRsFLnyoNJrJzAm1mJi504lCj8wnHkSgSJL7uFcTsSqNIwf126MVkWXx
KEuvrES3LdAqlegW2vrdwxnV/4KoNT+SyRRBT7v8JDhypJLceNauObP1W7RY0g2bY/QIcaU+bf8z
9sbTIWkCdO8xYCw5fQClF0n8T47q60JhsDya0yJ5xB8Y9E/wpOL1thpFefrLoHb4w2fu8mujdGvH
pGevD16svHxF77yqkpRTjCAbvnaqH6uquS7zu97nJRSr7ERtcUEYigWum9OGZNYa9CocZR1ote0I
IGht6GOJq6nQxlqMgaZw6rZm0htMqVit+qWBwgh75CnfzKbmD0cYyy++cdgfveOdUaRFI9Zhk7a8
0+5mh9ljG8dIdUZD+gs7PVHyodoOyPEs+AWtY/1aJf9UJ3chdFYbMjX4BKd4vfSOmeWUgkfZ54mN
jvgctbOa2zCx25bBMOnbQ8KzAH/tO+yBQ4/QqHwZ2Sj09w9bINvdE9GTMrPYgg9rLmsfgCnF7vtg
zqgo9TDKopZcW47MuICP0cO7ODRL53joLrjONQTBV6ZCp7DRgDhaCkbY5eqMzacCSvjZ/pCmpDR4
FuPFNRgLnL0pIrWIdsVv7tgJuH8UjcgDZzVA2INP9tLJ3JIKXKQX3wvMTIpRgSGEqcHcewJexvrG
Gsk5ofSWQ7E96DSNyR2wPuXk2eAHCRmdOLC7dQ7O8UzSdNTZvxisnMCQXldHhUURzj4fmFtr/M7M
8Y7DqnXHY9jU4dlhJOix5dbu3DBuFt/dgQz7WHP2YpKOlDEPl8N5x2v3D+2VVCnL/CGN1+IJqF8q
mUy8tmuhUjUesRB9D8yIj6D/h7KpzSZelgiDkezniP17G11icImrruuOi2m5CeNyZ86EWvBXsa0E
v9XVojDBBLpyahMlXbPyypGtW7RbinNITHMf1MrS+g3z3eGoKAB7NqgzBUAbH/7iOMzIpAsFJPpf
pGrvY3vDXulROYn5G1HBVJ9Z9w+qwNY+jHgg1Hzs5Q0gj+K8xnneX87jEizTV/I3EInuHpqXkxTO
CtrdqE31RabTMPyqEzh6vu/ttdl/ZP1HDuMXJdS0w6cBnfU7ncOBUbU9ExpZSSqqkNhFtQu+Hevh
lqL62+zj+BjsgtPPMvVctcXHjENOYbqmjB5UYgAVmkyuB+sll8i/zEoziCXyU82AQUgsjmuI8akt
1a3kZDY4uZgTCwkc8yjB+vTXObYaKDVWPbPLYj+1VAx7gja06N/BYGcrn9kGzlxrqsgvc3/TBrs6
HhfHQVMVlO1wgPPWKDgjCgalr9dO6k9i0/XdazR4XL4fH/JdH5z3+nxnjWcedH9LFXQbmi3DIl1m
txI8EZ0Um+QfwITMYJMcQK3FvSyqLrFLJ29X0PEM9sI/+C7N5mhkn+21qMhJzwdmqUJNQOdcAEX/
Mt2O3s/5psa1pVVeD6nEGldWJ1dLgRP8g/T/LlhbT8+icMeeiSr+Ln1Bz80PRg957ueiCTpLuI/D
AovBa/u5GDnviwXDC4A0SC4iO4CqgTh3/iVtscaEOB6sD7cDprjZb98LtfC8VPoWXuUtSEN8Pq6q
oA8e3BDu7o/SIAHUg8qZch9C4xBhB1Sju0JLDC6uGSJt/58I3453dejzqyemva6cgOBJMV2EnZf4
Kv51YiJ/wA3ed9GM1l/3ncb2bfdYr9F1e7AuWAwpJ0fFdwwsLHAqgVqHeoT2hKlwC5DaDSQQGSaB
Inz3RardZrC+thovONpGTLj9LUvzGLpG8jl88DGW64M98duFOW9Y89F+JL9GpCyD23mpTA28WMVt
VtlnLKsCNsfj4cANw1YL80lS6dNBtqlEnfq+wDxeVsNXTHGBY0MlrqR4foACvmnn+NbFHOZgcZ/d
MEOSN1R5BUe0y8CGvw/M7470CPmFykQDsNaICDnknEjEYDIkRCav7GJL8wZWo3jTHhu74SAXhtRj
l/l9uzCfW6cBZvNI4F9EDXkorYXeUfLzx3nGoxIHk8+NIBIl3K+S6W1vpJsqPslWMEWUPpbTll5U
LJGg1YhtnMxScs7hVobqJ+ZTFM8t2WT3TojDiAqjY/2GZSHJD6wXrTQaHIWcu/VPYF8Afrc0IjqU
DMmsi/0Jqa5e/tz3wMtj0mcQA+VBguK5/u7sYhDsp+V18tzHvrfGww9E/tdJf1bi+TU8IU/DbnQ1
P77+a2ar/H16hGWVI08SJ9CbNyCjQN7XX+KpTsXkGrmzjSexfrtVXMDPqBn8Y/dG6/YKcbz0W/JN
BfU+IlTW9enfJyfZBbhDm3dKbBBJ1LvUCli93eiMfOI5ZVobI+/r8Aol7bm6xIfSxvEdKV61nxCt
UPyOwzpv+v2T/LhvnQKTiAyclgPZVCu7BYazkf2Hta3qNZqPfeU/Z4DyTT/91X0MiD2tMb6Z+3Ph
cWcbY5iZn02tsiRdCmFFrHwHqzVc0RtfOivIOyqimimNsVnGDBxHjy1XCdDMCZnQSXAii7IAvuPw
AUpI/oVHF9QEPZnqNUJOUvmZ17Oajq8V+GXBCLfNzZOvOCksvjYzxJ+ZskQrDSHTs2DmsdXEdfgW
GuNxOlQ5SaeOSfEY+fgiJVQtGFTEJ/OxBLSv1lFRpH+AROTPY2ZAJtD3sB4xuXFT7akwN9FlDDsK
Y+F8wHCD1Qxg6DU8rVa7XjZFTfitfoonFfuVypchPwvArVyNAqhtqM2fNs0VZ2PIjsHqsTHAHw7Y
U1SZCmJr6oj6P6zbFyslAkjAAxaFwrmnWxgEErjrjvLCSZsa8hSBMjUc4+2yxUBAFbHYdDanmNCP
1aCAmBbaaD8aa9f3FQFoMRBq6XYhdx3OoT/BEiTCMvzYhHtyoiMHMygU4Z+9Vc87zDEZikIoyi/f
33ZzKUPnz2Uz88erTASIH5LMCfXAKxthyxjpNu/bJVLIRuXdX2x9ypS9skPbL/J0ZczYswONqqCC
hKsH5SQHNShW3HLKL8GV62fHxGUSOhJEWQEWuqBRd3m93MFJjAsj2vceeHRHI0RESlyGCudB3/bt
WGyeigiDw+vzN3UlHOi/oIS5w5LTNdPb8xO/oLCEtA0KdterBdMD46leThVm6n5txXqPBReu0YTD
eAZ3nCuq0yTSi5fraul+nvwMEVDhLOQO/WIBC2YcpmszfSe9mIn9Amh0/iZpc0tUOFmzpTGWsIH6
5yjuhGLVsEpHP9NItliHQg7bXJKTZkDKD+2uYQFN/gg1kJ87DmAPN9i50smP60mOu5V7Fv5uEMQv
wjL9AnDbsw1vbKr/5sUqV5VTVAHLHlzIDPxPOJP+TLWaP9OjYQD+GahkkKKWKkRkrsz7y3ehAJH8
6ebtXsF49iMhS4+d3Zxze0jMNeuRDw5oLhCDws0D+uK2PqcYkkx7c1gfIsEXGZSpYGQ8UFmmIUkL
uBhPo/riq7V2UGoR19Z9gCA082raABd4Kvb/8j/hVJVSYAbPZ8oJxJ5kXDF5EEd3URgeJ0J/Mli9
JvzvHiAZDYUDcqJ9HHTSZjdc9MJS2myepT+ezPaesEXNO8sWdSdfn7qVBjEByx5pzHgQ92QHlu8I
bAsLH2gmVpz/S3bh4FNla1Ax0SOIBizYRKta2NtyuU3X9YmBZ2vd3XQT5ZfpyyB4pFqew1CUjxoW
ReBvSQuMpN54QnAZf28J44y/Mz/XxYlqt/BLTs7bDoruammcQhBI0D7n+GgxDtPiT5xDttIvy6dr
yvLCAL/IY32sCyzuOhnm+QImuOmW8ZLQ0Xc2bX30+/p8g/pn2KMXCdEvayn8bXCZ5FWeWjfoThph
W6C7Bi/6ffgCY8X6q3swWCuEXw/y0Lx4iORs28FVt+l1LOWTvLu0ZVdrXQxN4pePOo/dhT+Mwth4
1TvNG8VZm/puekDRMk76byE4z7bWKUXFDZ46cYjAZ7XQk9/8zkxs1uKiiQtLr1KbEBrtYOTda6j1
a/p7gOxc1XLVuxYf7LpIp2nfOygk21CMY/dQuQOa1BnxmtWQzF5hh5/COcnIkUAHJfChljoLIbds
dwbUkRyOKUb8kPsn6y6MPiDqJC+U+O6pYs415YTsBAsR7wV4eUNrRsDTv+DD96gNW53cfd0xshhm
B8OoPkx77VB3lxOXmUDMb+9uqgZYUM2vpEiGbqPxvSvWFCjWt0QAggKMPy1c7QApftjQUt8aKtcZ
iQDBbGPfvCFCgxbNTsxlIuAo1OYmWHKrss1dGgChPrZtDFY7mPw/xy4iC8UixNp+DyqPeAA4+HXj
zISJXQD/uK3NLrnDngpwjYW9dH7LzCAN8XtyzjnifI6RMEqSEGk/hcPtlFmggFlXKvrVjwvWuqmw
Po/fYSSkn/yCa4vlSp0IGjp3pf7kt2rTBO56xGDEvE2RYtahzkdiVAIavvOsHkg6+OELyET8KwVh
Hmhw9CmdqruKaDynfMziaEJotilJOyFHEJmsEVdHW9bsVdSX8gSq0r3ibSy6gCJyQ8PzmonJunTj
YyBg4BgGg0OsD6Sl5qxwrlzx1KPskf47Ino7VAae6DVxuTnohutBiR6nbRzDWqce9X3QTfivDAuv
WT7y5rI1Oytn/5j7dL5yD63EGD+euX0y4WJZrQnxzLGZoo2j/tKXTEHqEwlXdDBnTieujVRayRDp
KD8hxOwICMIzGM8wHsijnkRZJtIpO+tQxk0bwbUReKVyhOAo
`pragma protect end_protected
