// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:33 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
buK7Lk4Je4KbU/jTqelMV1BRF6IjBXHi3QMxe9r3pLPClqvXsAqDSoIb9/A3PHOB
EDnXkKvi5fg+lR0G3iSJfI8+5u0OoVeb4pTorXqd8cVkPlpJTnddbYPGICfUo1J4
x+w94PfHcVvMWkbBIiLI8BTdB5gVI1FwVMwyFKlLxCI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3040)
HDJQYZlKzC8WDd+mpoPQfzldp+XAOykBaFKlRIgug8cQnA9Mz30Cw02UY/ScZTjy
kobEe5BOSxMPnQ4hqq2/+qGwaLYVaUHCpKk/VnbQTH0chxNhxYKPN2IM8zepcEEX
upIRpLYx14okwEWITyVKmUaLwEZ/fntI0tLCZXfWepLczue8heUNKhgovrNvyH9C
jNsTm8FdeKnWqWsAvvB17zJhnkQNXLezm/ZTaRQ7KYPreYxO9nH6SFVWgszjQ/wy
3Nla7P5JhXzSuFpvamp7BXtXO2WpG4S/Rm8MRY3MqmWLZ+PmRt00Py+hDtl1X1lP
uM3ZqWvLVDXJsFaBmHqGNIDgoQl7GMBiqrcoMIuBko3dj/y4vz4CPV2SIMTHGrov
qoRmsEmirrXt1PX/ye9x++onoH4/XwQeV+6pznDkTrrkrSUm175OSY6APRArM6XA
/K4pg36WPSsNp1k5iA3C7lkj5Us+XUJR/Bo9RdbbBVTE5bvyGV/tuDOi+6oj6FuS
FVP9XVbAO4qrGy8DYvmEIaSPiu+Nhu9p/aKDZ0r/Jx2EWdnIjiu7ULQvvrT9RgJd
ahdj3Tzlj0fMEOcSed9AAA6b1Fo4n9IjBMH0asrtp2EcAZKiFPP0oM94qMgLiRBu
6VsuMIHD+nienQ6jqXw4wB10oOGyRdkO/6TIWXtAC1qMfPQlgBtgYxN2JuDR3Mmq
2L9YX4shmvafxiHAvnyor/DlcGIG6cEjV8wxIZt52M+J2fcNGryw+fkDAfwziRni
NnZXOTQkdO04KkactUx9jfOBBjgQ/RZcjQk4QRLvCVDcuGal/TO+gE3GjTZG4dPJ
LoNw0d2CsMBGFzNApVsNWlzGuI0jPOgJs5QpeBuBDMPd8VFF2b7qiCRrzxqZIL0P
u8FTXTq46ngzEP865mLIS8zBGUpO1p5mRBUaD1gaWg153dQWNEurc0IcFYrLB3Fb
m9yo8qIPnqRahcRQYBwwYin5+z/NzUWS3rOW2AljDUygs3FdQEHJrrq1zmGM3lZV
UQyY7S/EWNDbuIAkYUgy0+CYHKsIfxyoZ5A5B6fHomzmpwCRfH/22JJIGihJvq6P
NRoq1a8tybUUi/FAcgnuLOwIwgn3dnherq+nSHyRBV0eAz1Zj+zZnuiLk9FC2MzI
2gOmHEE6NKc38S0t8c1e21e5ElXHgTLBdX45385VEGuYT5sH3zH/4DqiiznY4BMK
N3zEBBKeuRUabTp9Yqq+eer7EsnLcjnUf9R+/VAgn59wyxeMJDu82d2l7sUoGqqJ
VW1ICLlnK6kNXrSkh/78kqVQJKLg9ZbniudxuAcouEiDuLLRpNWQJ2vFEYxF9Trc
Pfuh7o7oYvsVsq5MCZpQf4KMKFHMLK6FcWyw6WHrg9xgZs8dB/3ybOzqd83adUZ8
2F6Jfw8LJHYmPLA0ySBn868yhxlDu/LSVDFHObBGlXPxiXZ1wALVQC1gXnCzgGeq
VGVnzZbna8n+9/EazhUNvEaXi7LQ8q4nujAmQjGw2D8NTya1AsDqZcE9vgEasYby
ZZEVKi6hn2HMIuUvf2MrJJmelcM5RZspMfo1aBmg2D4j18yBW70wIPgE+cUmqc0R
OsBspcF7OOfcxE90/h8ldBCHkMJI4P95UQNw51z6P8eDgE5jTxxxKV+zPW/QZgHd
b3srrFeLEz8giaRbZbRYqyFpw4pvKPUqXa3hDjjPG/ky9V5MrBSyGdm44WGXwrlB
kPj0VAZZWjyTfoYlBmv6Tc+AsWmvQVK7fZ+XD1HwyhOn9LVLD+goAzNvNrX3Da7s
oYQT080I2Xz7Uskktb3CRfZEe5FKCyvndmaLsUPvRGiBcxiKcneVA+byhmfcQUAh
WrotHQVlYn7IaYSR5adAxzTUd+ytO5xA8a6INm6cTGChpDoL0hzCJxFXU0zCDtvs
arfUh5ZlLTYzyKZQkaKAd7UeCAW4t+hijOmZz3E0H0jYz64jPBt5XEXTIf1gecID
/H4ZuImqLjoNlFNRslbfceqoIqeaIk/imZmxB5MMm0pmlzEteSXPafZysCqZCN1b
kKzEdRPItWC+LCKTOixkqTKHmp+hFfb1oDtKv1SmHM6lgiJOHaZux2Prof0/aCKj
E0DY1O9lbHTVJvddpnW5drIpFV1y4zX3OhzHfW9nwAW7LGTEBDh/VTAdEnO+G0kI
/NSwEgsIU0LAMO8lk/dMpR9p3EKPPD2boxiUpqOmMnyWmvadBP8cZV6OpXGhiceI
OxXLdMNVfPriBo9nFBUflaVCIJBF+StCw21xUOTPxlcmzT3qVnf0xR+h1ly7220M
e9nFYBeWVt/kSfLY6Xlaowjtr5J2c9nd3L3p9E5Y2Q8yA2/yTGmF7DTLWRH76atQ
eEHf9hL+hGw5x9ZKdDvOIx6Zb1p1Juf2snhf4vlmQ8QRiZ5fNor9QMTZIIMHNUr5
H+XbTtu2aNiHFHCiPye3SbeM6QqLHN/UMZwRW/lZZXyqzHrR83uywlhu9xcs8X9J
D96z9kq3RmDFM6N0OZwGDQB6UxzuPxu3bnOjNs+VfbAx7pSDIan49GzxQBWgVdlU
bUEAyMe7PZbs+cpQ6DMmLUTyHrBsAKNXTYiQLp0OPcZDTci50gDORidUE7vGb10j
giwpCv0GlGbpYZq1ol2UhQEYXQdb+eUuBhCDMQPbxTZb9Z0anbsdEl9VxzhFoB0E
wavRpebaNH39A8yuNEpCCrr0OkrGFCr0/aP9z4OvsADAzMM9RReAPtPKbnQapNxZ
Qw55bowfj/iZJDzTreFWOFsubUPYwMlnF+sVFDqIYf4K7YqhSKSBEuL1Ogi/BXSu
Ry4c8DD8THJ7/7nbCl8UVJzljt4rLOTrdwwm7W9mrqd8Uip1DJN3kEw8F5fH4yUz
YLn6O4+r5FJzjMXyUGJlj125f6XfFLi8oijNtYjmaWj6f3uHfh32yCqdtXHqSjYd
hHJF15Tso8FOUGsWajn/6nbsTRFNv+SwvT+yzRTGLDQf4kyqnrdkCtj0FfRl8UjS
5NDJCE6Q7miSj/4UkjvsloLjHifwTojliGfDT5uEwhkPUiPs5Ht03rKCioJsON/0
N9zpi5b2Gkdz9Rem4zD6QX+FwMwnyftmy0BZEsbiQj1Lp9TSBEXAJHTtRUkyOSNT
p7C4/yrxepg1SbhzfEXVIMAC+6a71nhnoqvl3/q87PtVh+nwoe6JuhiDhbVchczi
x9HhgQCXmrLkufZ1bpkYtUcUsg4Ayi6kODK2UUT91d5LcoSl/iXlLdq3Mz/AIk1i
mi8Io/JeNRzUiqiKbjURrsx7H3YemRqDlf7ptGyNvBWo7oYo0OVEm0nfTiJDfLvA
ljoqN+9rTFcPOv9iLEchoj19g0dA+BJvuPz7SZJbcqkwgbuJCTaPigurufAJnyWA
LxpTV0VRwogxaXFktEpnN7NGQEBaXvvoaoO0f8ESfV73yza2CpC6U0aNXqPpWSvL
na61bbbY9KO+o6zD9g0lCpZeFTz2nU4OC81APt+6RJOl9OfqHvteVdHfpN6cnQoP
B62CLLdUlM2tW4CPC5iYbl+ZY85vWFeDpsNKxoz/nI63IxZ1NmWFdEM3g1WVVKdT
SILtwwgg0WPzVx7GbPKLo8X+4YVUIWmwI2oDOw0xANxJeuS2f6+9eRcX2ghncxTT
i/Q/iboFYNmK5WtfaskX0SLTTNqJFwaJa2UdYMHXibiUJ55bjwKnXX4HkDGVX1AG
CQVX0DE9wTRWmWk35wZwEd4aJ0oD6FsSEKcVFTJSTZr/UcKclSAICx1VOnfrpNMx
/Sng2Wc322jh2vt2JXMbbd02uBiSloh/U5bEFpFXkMjsB/FV+6htbfVLYIbGzsqG
Ajg5rNF/mgP78JU+4pte+jlvxIQKd3oJrbhlg07yWzehe4S55BvSBGgwqp/wId/5
WrYD2MOZHyEA8r6u9D2fjcZuWOkMS3TUXInBOLsswyAWr6ZAZLLQD7AkhcqaIKZg
N2ZqLkhzB2cOoi8Vrk4QHNe9M4wec0YCehGskiRAt+yqcEON+yQ7vn02Uq5WdDx5
lQbfaQoT077F9TMol8b6vw==
`pragma protect end_protected
