-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oJaAgHDYTVRiPPX4UiFq5rp+emp78AYvAvGRYfyy7OC8FIpNJ0MyzrFGuBmNr1vMJd4aoeUlEBgb
5s5uDyOGUuBFr/Gyt6Ig9E54jn+7xJy+X93O/q9nJQ1l3vUKYbpcmcYOAb8FYEN1RRnIvin7Wy54
643F4FTqO30HoRIt2QOGW3TiIKQhtbNcbSdeMrCwjgrT1+fItMW1IyrqpbFLCkSTfSkK+ObXq7Rr
1kMWqUr5QOk5/GWFMV+otte+AH24gkT3rB8a3Il6XZbjeTzQRd6L1SkzxP2fljv115PqNg25mOvb
RiszuESpr2JLCjW+x19HliCIdtOeS9dXPTlgaQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7696)
`protect data_block
AkXcNv5ZrxeCIJ4u9sA8zkEP5wWq72U8F7+K9ZZ+97BL6TFX5vH10Y+1b0Z8B1acpITb9K66NzO7
glopWKYEJi3Ewhu491a5ZJoWFsVRaVU//k1ek3ljdXfBOOHB5fSVy1NmWlI+9czaorSstsiz9f5i
igtKROxM8mObVOL8vXHkFOKaeBzql1zX/ymIB5rBM9+PC/g9PRYWY/pGyzd4dXirHHBaHnXvQTxe
vhqpL1jtvjS5npiMtjcsW51P31YMIi4pS47BO62gWQt8L0Ku51zrvDoueF0952MuH0WEe9XaO09o
vz71tul7vvO+40GlXwwAci3dfYTuEi4EBY4DZwHTwcLSAwllRWU0yRJ8863AJndZwAq96v+YOH6y
fIXtv2xOLJqjAQZvMhFBZiNviEckqGSDBj2omIBUj6lLydlCzz3rhiD96w0IH5nVhL4CMjtiZwWu
NsrznzhwPEzfvq8kCAfIlEFEpz8lDYeVzx4YUwAYTBYZBUukk9LvUi1h9YpB8x/1lpyy7jy0+zD8
BU+0Iip7CmV5n7/CAm8Qc5epzPvQDktl62YQ3NW0FeVg6tw18+8gR/YBTVLngQTRIbw2f55VLYR3
zJ1JNxNff9rKJuSiWgu/WELdJ/4a1KvGAGSxAPxqwvItpt/Gj+rPKEoHAI1ZfwRwclQbkuZDV2kY
ejt2LilKZqPvCsIfdYvZanwssmO8/oDRh+PJtw0C0fr0vhTpV8PT0jiJCq4iPnzs9Ab1r59bobjU
Kuw4E1TavaKjJRY6LKHeiSX5BMSWNHlfHBvHSwZtBO4HL/oVNT69hRPNHLRucHR4dphzhf0VbL7c
yp72qXKr3+Y6viR02vpkLbvo3ZE5kvQBnVKyK+wH8jqTLsmWREjsL/FBkL11gZgAJPf9tqzNiYfe
exjT6CxHWrmNkvp9Dj01cMGik0Ah59zWmhrr2meBm+cNmAtzsEsjdQaFi1Mp0XhgDZfLO6RtlNQU
1BV22b69pg0h0gRQU3e2tad5wwV21CPsHQzNyLM4QKawbeQEjN98oHISGQUgazZA8T1Hpl3k/lMi
c3Y4kOim5mxrsullLyTfqvFC1iPz6zbdnwTnYV02H8h32DN2XoaHgSN33eo3Vixc5tN84EqQ4SZe
OktL1SSokef9NU//q+I94P5lsL2LjCByhSqp7Cvd9SrdDctUeFw9wcc4M2BAmYjOJocjIiLtzRuN
ylO8sSvAv1X9WX8pZHrLjuYewDmPY4PFzepkIifath9mBMoUTAJfkCzEPViHgQAAKGvsMmv676co
RHmHDdhSt2UNr1SIw4RLjh5mnUoxyk4q9aDETWVTyqNnOgvHyOM/o9JSBh3VbWhRX6dCLnaROkWl
q2K5pnzBXkZgeSkBHZk/QfwzO1quHN/YKH60m76qvNClHnNB+g9K7/2vOdmZsjjxYH/42jZVcIQ5
JAPbicLwbT2YByFvDD1unHlnQoZO6CuURzFKuDkWvVyXnF7PfnFnx+YVeeP3BklJutxM+lR8kSLl
ESeTZ1w9x0lonVn+gTHeJa3xSGwq40i4upb5agt45chXmPLAiTTxb4oT+MEs2c5tVrxFwTtD005t
9c7omqXIApPUG+qL4EraZTwBuZ8vutKl7dzDHTCmXyg7KBv4TjY3nea1UYxpsC7AZG2S8VDLjqIf
2VJM4l6NzK/Svet3a7pIQ1Y2mlbbZvctp6htq4he0MfFyv+R/U8FCYW+zmakCqP90O8d/PKy9NYc
oXtAT9D5J5EHY20zcWvJRivogIgw+7r4Sqyas+FXpG3A+S+cvNYidv0foZ7+c0MSNdvqOYfXS1e+
+D62vH4gkAWWQoqyty1ww8VuADQ3O8kZ/ulmIslNKNeYIHpH2XfMJLHxLJkKt3IuJ1hkSqWoPzTr
XXhBBC4uFY1s30WSZ/R2Wmtf6HJeKrY03+4z9+gcZJn99uQfX1mWPC527UIl8uCYwUqTg6F2g32d
RvU8An+erlmA6d9Wmbu3+A0rhl8Krem5ZkkIQLzOPza3pPCNSkbwrINRzgk5eO3YvTbJtK+QB5O3
Vplxab8YUVXtjFpBO3WTiL/zsJKBnxDlz6o4ls+gg1CLk+rHDbcjhu8ZqaTOECtuwfuVGA8+gtdw
m2bHK/hQH9+sq/VV4EeMaGMFmw5KOqBk/wQdWWU9bafBeWB/CKSQ7cG/7o9lgE53UYsJrMYgo94a
SAyj5bDAtsFPXPC66TCzdR0ckOAAoeEnUkei6+bDEPHTfS/CUE6R8ohrpfO1v9tHBgdZ9ZNbAx3w
6LKbeLWNvQqb/lNxXV5TkEzC8a4fnV9ExOk2MH/oZ6fUzdZJfvY3Ik7NQCND8hcWA/onjT41tJW3
KMmpWdzhb5PVMXZRm6D3UzcQqtKEQgUaQjYPL6R9bvibVYUhiYRwi36qZQUvMCgUxSm7l5wEFOVh
NnMA95wSeqL/Lo/asxrVaFraM3K6Fykc+hXYizZIE8mEzDVlA02ZhYlwmh673izskprINFqbQCar
brqk9lCwIOF36Gnnfblxx8to8IIl0t8CYsavhK+vB3upYSoH59hnANcn7XfQBhfqaChBa+8LDUH1
rZLJ0TbXthjPQ738qXLAsLVNs3UkUQzXWqT4fwoTOh6LlAGF6xOMxzspPQmlki15TZsP8DuTn89a
UVrR8ie2BFwywNnou0mLAJDuJDx4Qg5cTnaroqPk+UU91hL8qlnxKpGPw6iWkEipYbQbDKHOCkZK
B+ttTH3H+6H7Ilfuj1TDo+13EXcnZbeXtETQsRh03VtojofIlrj2HoOs7Hq2jZhtYKThtRrVCLBs
IUFg8ZePwP2uHZ45mIHdeoGFceTZwkikYQAg0AllbiO2Vjy+NeqgnZhsJAhyV01Kc1Fsjck4lm/n
VBbYALPcovC4EQaljjcenN2hWhe4A3MO4VsJZcF67nalMFswHgNqSZaNxnEdsl7zIP0LM6ZPBteg
SynymL/5Oy9M1Rr/WLGs67qO0pnEvQz6p6V0qsHaDxfpqkCRZS2QIKO3IfF9+jGTMl2sPJzur2Ze
4KxUumo/zk4pLTvaPcAErlb5pVV05f2jw65rZLEVWJZ9A4sASCx+b6VZHo3DgkYYPFmLAS/QoED2
aDP4kaR7SDE2APuZNZfDP5VqXYJ/fNlAWCQhAWlKOMKrs4hNfp6e6Rso/BOuSw0W6DjFp3pHT804
K48fAakdP6U8ZpQG9y4YrDVXzQ82dPUYV3eHhKFC4JxL6oM7+j4h6g2yWqvfby7ZaAtM1cAAbB8Z
DWd7lqBjex6qj1YuNgWSQQgNJOgyr99mzJUVny7WwfwBRGdkziRljNEopYKpOnl/dBEpIxMbNCHw
31WZja6iVXMsbpoML3Tq/mEi5QlS3CeSV5lV0BxgkNesTGiDyaxtcp0v+MdH1pqYmP+VIep7ED2P
hjXTQn09HjZjVLEAOm+fzXWHGG9B3wmXIQUhAnzyoSAvb8AqrclI7Mjp68fWe7IooowHw/qDGHIT
oHhS7Mv42TC0B11gYWJ7L4Ex6YPw8bC6UmBcJPXRPbrzufYtuWuugk5Q0S6gvW6zmzt+INfW3Xb0
pMiCT8H20t4+DhO9E1+6ojPgC5JpCSZ2qxuCb8vxqMZ1/4G3L+ibFAwEHhpqDiz/gXuHzULzesWW
27WMv3V48bBEt/5Po6zi6LR/hS2Uru9th6OulAT/O6SlS3rIGOQChfLbvqshz3PSXBqlgphxAdT0
F2kPS1pWhoinn4QAJeTjYkesvifr5Jv8A67PX+gPEyW+alBQUn55RLtCnU3Z8z5ahU+JIJwTX3YL
566CuQAl6PYfp7zyHtiRNf8vvGg17CQCYmIbQEghuxs5qeewJJ2MgN9I0Thi02St7ckoO53PCDLi
GHBLki37nxc9JKd/9S6cmvAt8XLI9quwaR40WX5yiDVcl9ZYUP+K/oaLuuQsVILI+SDoQe2GvDvN
SlaPSF2AQJAhEe5I/wtfaYgK/J0Ctf+iTK3pblNp9iBnaYwcI4/6E0NWXPL4yrKktwduK3W8jX4U
JHPwlIGJNsQgaugKV7zKaYFPkJixJqjk1OF9QfDyJpOCm9czdIWE2myPQBhC93p6lYKrxvYjVSlt
OOgwwFbI4BsfIU0wwVN5SBK2N78kKzyxzArgUNhFHfbUPgFKEWtgVmTqEHJiU8X0uPD9Bf35QZrL
FJdad4IZYYqNbZndlpQuBeGfPlBjPA2MRE2apTaEaHdwypXTs/0/vv40EvBr/b5IPOih5xZxxkWZ
+Noh1zFkLgN4DMPu95zcGpLGWOmSWfnp2Q68a/DsSVYK1PXLxFNq/ihbT0XDSaWPQyxl1zgWDeAO
+QKKyLICa+8YswNZTgWrGyrSucydJru1LLMDy3mNbSfk7uI44I8mFBVI0CSU82vdZ08ew+PtUWzt
9UfeUoyOhCLPGYm+Fsf20MP/XLDafXTpnahOlqCZ9AqjlLO1hkMlwzNQIstzVMUsunTgjHU5vQ65
Kr8IUVRB0IMuxWcqPUqgyNqTOJMRLkmw8yrglXlJncwbxQ4V9CSXpBaTh2qTrLhLhQTodPhqhc/O
+I+s/i6QOUTvpZ+HHPMrDxJbDbzNknq6sqRGDai82W0ZRyHdRKKbcjAWART4NMY8Kjk2h+1psiNl
vvqnp1HgStbgutZV7GVRsgOCEyrJLeMDc/vqmoUWV5muFl6OhRpO2XuVfgv2+QTJKd/e/ccPXgG9
zVzfdqJx+A9yTiGpn1Upjt6Y1MxUm0GCQ96QUwLhlM0Vj2p0Tgvz73naBHLAwM+0GWlnrdD7SzbQ
FFPUPTFnIw6Rc/SHO7BsxbaWFrs7BtL2XVFwaLGhUmQzwLle0kGUUAZijXgLbz4KVipBa8DnuzlU
Dt82NaNs162sSuS61ULHUGQiUTZLWciziUl+Gs6FEHyWQEKk3T57fg86V1GP2LuPkzE/vP67n79g
vIRjN4vBlrQpHN1LsUtQtZkDfq5wUyjn5fW2pPGLitb8os8YsTDMwSbVH8f/S36i/2sRzKM5LIoi
/iY611Vm9Xbv0SG6MJXeVp1u9ynV/MtTnodJeMZapqt2A/rDiDzylc9dWGTKo53ejnMHiR6I4U1A
XkVvOUIN4KGP9ahOXdUqm9Nc8JY17ibg1E970siKQkvlziJW/LBL7loRGFhaZODqHx4YptEUlDXO
Wg4CDZWNZeV62pB8Hcv0G8MtuxIUUTOo23vxDQ/FzSPqF3q3PpFHwIS5RbJLK/DUXr6oixWWpBvy
IKmc9PnDedt4dJhQD6I+UTuuiUf81h9AtEvWu5djG/xCXkHZoOEL87Pw4QoaWfHGIsullb7m21Bc
UnQ4ZLIsv3wClVYgGG2yCpsIIswbsKmimGTzeUkxYKExsxWZJYOoeaIuN6oCDnywK45fS0N9Jvv0
EyqwxFkspAEHMHI2pNCEW3GmaznnC5mq5lKqZCY0g5VJoAGhjzt13zPHaUr91SoxSub/3razEw5+
WqDrCwJF2xHqoMh26Y8cm2iDhZFkdAxAZjZtt3M11Kiu8X8HHB64L/zZV8tWRTzjaJUyVfwNuXEO
fSnmKz/LyuxcwxUpS5jHb1ZUF/kCzY8aDoxIL+nb6futz9M5+mV2VgZybuRP4H7maUcrWVUL1+/Z
Y42G5Zf0oQBYhCQMf0103KvOezvQ7JHsEFhjJdqi6E/ue71ssriSYksp9Sz4xZuI0MslrZ3mcfiv
Fqp5SbRMThTS47/SLiQuIITJ/6XiiiDsIH81CQQJ6AqJ/bsXdt00vacbXJBh+OvsDpweUMKmXz+2
Kf7/0Seuwyp4TdNWivCQoyqsrOPObQtzFykJXYkq6PdrN5+EKnd9Lyd+QG4D5Q7QvCP3hwCqUGxs
VIrfX8WlwvySpYRQpiPEjuqUDejnhHKvGledAYV3C6sOlFVKITBYRcrbMSM+s5PeMPVhjneJjdz2
SEuR69xhW0EnTmO6B6Hq3OL3G0k4lhPhkpKqG8Prk8MP00k75rG9ri/SfO8J60reYat1mtdrHrYy
OEdGkciF/LXULtcZieHwhkpAsgPWQ3DwlrS62XVXSiprPNrljor8Xc2t/ujJrq7c+EOSHkDwWXOs
/8f85I+br/1dmAmGPDgQq0R8daSqeJimZ/fL6333h7JQX9BvVGtbWpDEt+T3TXJBPJRif/xSDsKp
62Gm8VIAYELgA7RKow9VVHh4KLk2Z/NB4sT1XPrJcd0IdQ/FrwAu3oA6UwOVjDym83va5I1D2WJ1
qQizJGqaK/793yG87EQUam0FlwrZ60xJOR4IddRSc+5dIomTmDXhBo1Z1r1P2wKqhsOX9UvLv9Xg
NqYfU/4QCxb3Ie9LdtIFHd8WXS2ZmxEph9nhqVdD080uMFZqDoyYW7dl2u2NtdIEsWFEeDVx3fKR
h3CbdnOJbiK1oRCWQJnwpXa4x4ToTaaSQ4X0Mz3xy969rqnNcY4/Db/Oz+MqBISb8dvtbBU+oJaZ
ilLSL9KMCQ6+hUulSjR9P7pIEldaLO/2Cg/THqiZe/Drbvo+16LTA4c0RgFtlBeYVZot/0L6K2PY
mwzHC44q/P7xHRojwBC2rKB9J9pTVZARfFrPf1bzIKRX+ydtriQHtOeMgXCo/5OQKvuZGnJDkCIr
qO8lD3+lss93INLYjHhy5JDXJhLVE6sQeW5yI8JkpCrsjsoBveZogg9kbuGXjDfhdOYbmAPi8v4J
5SSrgX5msm6T6zBBab2PReDjX8H0dEUbcY6gd+pYzgoLEO1+Qv3o+4DClrMGSp52nD7snfQotwaI
vh+u3QuEwGuVvNTEEkZ3amKzF3MeJp7D36Quk3tzibojgOxIa0bX6Ex287NdueMLaI/g2+dFFDpA
ZLwgVwBevgiTdSvnE4iBDAlmubYOVUPTr7ibMKPlk1DuwYNWfATE4YvJ1+9GPmK2SQoZP0hXLHKn
lQofbVvY+deSID59+XoEIxh6A90BXky8/GxKAEFozGFZptverlk1Y7JmOHORYYFlpFistbtaic4d
xIPKmbRu7iS3FMwoNRupSO15vDCyguh3ZZGiwWcek9azJE+KvUNIAD2Ww5zIFl5lc0bKi3yEo/qF
yzlNO4Q3XjwfwD4oxlMnXe+pAKEZlcowHHGgiFMA3HuiRIz6wJ6gpm0+0jI67ue4nzkdg53bqnJZ
TYwjnmqRXvu0F+eSrDRWhQWmhkHhW9upe+IViR6Ll9DlJw7zHUmYiNABESMn8UsrzqnxElD6mgaU
LRGI+VtGwZKuMJOIEWDC2tsARAAahRNSWH5G3daUzRwNQR15DZhie9Ds7OKcB+EgJYuQ5/p1MGEC
FBtpgWNUQwJrJ0gGZdhzaNl3tHhRR8HGP1smhFPv46DqRcrA+QuTuen6FZURUtPyBv4OAnN4FPct
v8pR3HYKjcRAwVsCPg58VoiwQiAqDnrM5pq8fmFJyRgfThJj+qI02PbO29Qjwzt2yTW7NAQjFFUZ
2es1ZaRMCTJCrfOZSDLzcIEgCyhPEpY9kw85IXrG33dugM7U73YY6DMg1igtkxBQbFDl/Z3pXft2
peq1wGhhw2SACFowUyXFpVKCn+TpWrFsys4VSgXgrrDfmJRlM4PNZGWGGEsnqbBwE+hnpJPLfqW7
kA4kf40Q2+jABgjF5mEbLk3bepKXGuQLnkHMWlMcbL0TBkmR1iw8Tj40rc7OemujnlxjR74/xjEx
DBhuuakWF/Rt3QlJYMYqbub0wQBbAg+CNBbrFdc16t0JRDoTbA1ql1qztUrsHw0ef5pT/yRQHHIt
+OvVIMfATiU/o86sM69wa8JheTx56+TyBd/kIzo/ok2MeZ1UVCWc+hWj9QY4Cpr/UECxY4F9Qxmm
ofOptLd7k9Py5MqNURV4u9cy53l5qAXOOh6S/It29wUGF2WMI5cUr3drWiThScuwG4RBih1Va2go
H+uk6M+O0dn+ycgNcprXzUAWsHQUXN9VBrzj/V8CGxEVv+M3gtXDSIRYVroKQ82ehAgCiZIrat0K
y+jak0Ge7jArnpi9InA1eAsioI4Wk2qrDj4LSlL1jm4cLB9N6DsPxNvIsrVBZo6AqR4YRCD+rsX2
bNLU+xWqAmNCZ5kgopFMdk7Mw41EA8eNmdyK35wqu7ENOf4xNVSKzWO7SPTFFh5eXu7YqvH7vJ7k
FBrq2oQTEJ0Ydrut1vf4fNWmavaq8gSSG+pt+bhaK66HFl+dMu8yH8YUgSlQXwyriZoUnwbZeWo+
GjivL9GidiyDYQqPtqijwVraAPTk8AvSQfTXp35wh2NrcAkYWkr8z7+hLitmQwEe41TjoWFsleXG
20RYydvbbmWiA94+4IrLAIzKN5YqHYpf4ICKWTtZDMq9Zj/WoszyfVXnbO+wkucxgSa+UfkqYXFu
RDgTwI35kOvp1DVLQPF3AkhR4Ks+RtqN6t0E0xuSob1qGKmG2N86vWP/zxB9VMQkRRaN8tXLZxc+
p6OdPppWvIWm2UJUy7w/SiTJ2ST822MEWdrMZsFJOxVQNBXCWz7kOQpgDOjOi0t4I43WAXOYJ3ap
y6zT/itPPv4HYfQFHiJn/kWiTejsWyRL7kecx/AMvH3zeROxZyGqoB5NtiRLHraRrqvXVGUMoyir
12MFzg9M8aITFE+epG0hBRvUSLj6+v7HvkwmAy1LiaIKZXjarECrQBfZNae/5uScsNN1wS/1hFkX
AjmAONJ8fj9qrSqCAsBZTbbgi5VDiOXh8wWFRViFu2xGmcBfKBertuXlVBhN9gkzbE+lhy8X9f9e
UeNEPnuBcnCaKkaKWMMqQFNo8q9BQJBxHmycZ0rsE1fI3+xlsEQNNOFnBNKI7aWmV/HrISqfZE9a
0lprqs06A+HtfJmTW++VP0PIZFXCOr33TcJGhMOELWpD2VHR5IuuxVq2MCzd55C+aSlX4gfZSAYS
OpFEz58QHIb6QKek0goQ80mDo2TKjnKkGPE1kx3wEn30Tt5GMXg5Fx8w87PMHMnY7B2tznQjgdut
q5L3AbrPCwIS6vnCoOKWISW5wOh+1EWb354agJrSY0hRZttYQ1X+txGtFH91vNabXqGzeVBormdn
9NAzoIIlvBat4UcS1Hooe/wXp+IyDIx/TqluqUuZ637z7xMysZnvP2SHCo31fvd8sBsjbPR4IFJj
tLflczG3admz94NhcVWprifWiuWmF2Z1ylMghSONzZPpHbkLApt1HuXzoeqGcYEef7AG/HYwBsNC
b5PXWEqjLJXAk7/01N9e+PXNztbOrCmbywjYXL2qXbErCMpMUYjshYyJO7X978kvG+atyY40Ro6t
oPB/0dVGAVA1qW3NGRsYmy2FWZMNd5rLf4xdpmrOioobAkvcq8EtHyqeGSkqJO8IRTTqgOhO7jUp
AXx8aK0TTXU34+Jgatnb4M27KeIE9MDE3TgKQpPgZ7pG+bIXoRqHd2UHkSYFtV9taOmPREi0wJXv
VCzHvpJfkNBvGbR5jmHYViWkjPfB2ylnFublSVrJgxqqHfTvj5WEo3K+wVqf9lrZuyFPhSqC83xZ
zgF+ZU0ttrbcxdrSwW0mn1CI44hHDonRuqUBLJwX7MuLmYY1+PY7/X2hdagzOOrIGQPWX51A5Kjt
xy6n+n2q6tPKVXZJmcPPargehRL8Kp/lICtNvGjz4oCrAAnyNK7CMmx00cIeMKJkgCQ5gv5W7Ruu
lrvUCZlM+EUT5NCKtLnDDKn7l67nPvMeQ5/WnaIXxAcC5fRFaxbss1j1f6YBY9YIo0iAqELtzEQe
p9pwMQACTJzHFoeg/vZ3UJw6omw0e7FkI1wCtsZwjZd/mz5BxZUfp+l5vguC60nMUH5fMKJUJS8u
+FySQUcOOtvIRqWUGE3WagB6rRBwLvjf9letuiqsmzawXERBO2ac/3DFYc8Bn7syzMkaq/X+duzO
pvi9C5kumepG8lA8ISvG24c+xwQ8JsOPzDb0F4CHt3OkYoR3FahlQcw+E9y7yaOrsC9cP7+qS0dL
780Ltr0CsWkqG7V6MhmlZ0cnCJlEtHpkZzC6MLG7/+Z1AJkY3A63tmFlmI6rEshRcZkw2Nad/Cdx
lzMOIPSZSuoxiUXu/wvTjDqWdseEFDh0zWkaEjNhMa2xQAZrZIDEydq2y4d3I7ju0QANuBCPtPq7
vXkVNZIjkGOaeRzrd5zCZpOw94AW44sVy8WTjt6nSx9gdCEP+rMUMRkAF3HCwrJEbcHCCdnnXGW1
eXsBq3wp2K4/ZAytlatyNaLX5YYj8x3kl55nhx5c4yaWIqRC7M0h2Gf70q8xfOctOfPoU+N+d+AX
GA==
`protect end_protected
