// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:32 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wwix2r2QhbbJ/97YTtFSS/h4IA9yfVp+L29IsdfGU852vTjRCQZA7bpbc4JeMNEQ
xvlN1vgHXzOeAFFgy2r9jsdKbl110YdOSIDcVbICG5X6fDqMU0i/cYGbjtE1lAfR
lIrVckqrapfWUCVqY+MM5HWcPVXeT+TuPx7Ik5MT4rQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2064)
7eFW9EUxD3F26XK16KSgXTSPuh7cmWKD5MVhU+5owmUiwRVX/r9Vi0cvR49zLQrl
UvHbgHCXfXFybyJivyp8DTjUGKcy92fx+xxvTwVkKPUhNpOuD6xwIKSBK+Y7AYPF
81aClmhek+qag6hvSUfJ1uEZtVSByjqqxYj27LzDjOP7YZWN1GGRNTx4eiDuTD7f
ImbIzIV7KHCQSH7hkhMFFMmIUmfKmTmlztbiYsOgGvkOlpslBauSbfKgCizX66PG
YqBdOf7WzuAT35fGET4ckGkqzEab/CJUS1WFCF6zP9Wv4/Rt81LyStVBq4iCG6ig
wt5DHCfyx4WAZd4VTaZL1CW1OIYbmkQLtMksTzZDQFfUx0IwdP6EHsl61d6B4Uwz
BqCD+h5kyeRYTo4ADgUJERlrV2hUhoYSv7KRlJBhdwXEH/ztxoJV+BwlrgoN37Fp
DxDVN7oSTxiUKdypQwcWI7HsGlNmuh5/MyhQMVsnRLD5kAnZRawVfAe8l4TeNu8q
+3fuSMRPtMS1FMQ2KNCGf7Nh77jLx3003DekH5rqylAtCgeSZ7CWqmBwUMzpdZUL
e648ZlSa/OTuMZAvmkkYBAWyd7EqEJOvdcEamQWY059KGLeiNU6IXuCJ7uDL6oiQ
UfHcvqPllxAhAWgyAG2zThLEB+B1zTpB9q9rKgBpH3oxJpw+6SjGr7dvphvwoaje
5QtyBo+6AF79XtJrvpgCF5HklINDle7dVIhbsE+SlPqhUBVT+PD2K5kl6bSkgito
5NbEJvXSSOou09hYFFXBXModnnfyPHNXLvLz44AzdBYbZrcpE6u7O6KGKnqy2D4a
NFgIphE0qykVRQ897xvy3JJCURGoD1gU/wKBEUZJil5oXx71FY+VOUf/TO+uuxks
wwzcudWpgs7k9pjBBdG2HoIdtZH7B6VQzPOAX+iY2o/NkSMOi2cGCkCAnzrAMsF3
66UcdcT4KTxRmp6oTLIlA69E+O5pR+edKGJtzRydJdow7+Np0WFYbDIY7QrH/G6u
SUPr1A50egk8uF7BslRdcdDn5LmNFB68KQPWqR4ZLQVEzNlzObHg7rapGoDQSkYB
d4o7F+hv9Q4h5HwFVUFHacnBrUiGq81qsId9XNkmM1V90W+aR1KDfFMH9Pgy1l1V
D3no8IOfCbjmOgsscZ3VaQ3YKBdiJS695RX9GyMSFwEXBvwCm2fuoHzwBu6tRgOh
4UECZUNA7HolYEOQAhjNZ3y3qW9IuZ7BnETNFbc9AggoN1AITZZIIdPK3A4Okdfu
3ScYEXW/zvBOuZd23fIy5fRz8TAMF+kqjAhQ/oa0rTwnzZ5Q5HXpHSksVVQviKlh
BbZ+6oLqTT2h0QKCAjGdtTebIV64VETPckdan+F1hHQQLY3a8TXeSBWMujv/pgrA
ROW2a+KBVGkncQTyWZJ4wKkW6qTAtatEjztARZFCtQxscMsHONAX0Nb7osPal8L6
BXBZ70gf6KJtxKcgzOm8poABmvi+0N93cKs5mUNR7DkMaqHotGnj9VWlZDgK1bwP
pVwrXEYRM86SUgcEMpmMhIM3t5L24H2GUtg25nekYmQnzJGC3YSR8/RdpAEX8s7A
NCXutpAH8rtGe7oxzC6fNThnHM+kNwVJ1zGHnOSTBsUAZpOuOZU9bG0dnKitSEp7
4+GMtVVJpHsOAoXLrn0kHi/t8bWN+SiCmV8sEcVaPOqz4L5q+PAXT2NwihmSLm/J
RbADuNz4seJ0Ptg8Q4yUci2wkNHB9EuLQLX30eMCAQ2IyhTNPfTT/tSnSFGGDw+g
J1YQH6rkwFSFteEkJUxTJZ0oxb8LnYatwtPZ+xyv0MIGpgYa2wDkAR9mpwU2Z1QC
vUQvietxUZWpqxbuICyQS4+0e84f58cPhvq8GHMbURe1SXVFWHmdsyQJb03n9Ngs
8qBUgMyC12h9o6adTxs0IpPhh9eWoRZCfIlHSqa86894lqCOXsYpMa0V6FpyZC1Z
HoIwvx4u6XOEduzAatMMNcws35XUgbSaLmRn0v55W/SNvcaUng40fjqG3uSHO+SG
S6av0HyzZtA/TAr82TCZZCtvzEOVyXTCAFPDnfrHnGyN/qm2zfz7jqbYPu3irW5o
2HmCenfwNp3g7BOxHqP9GogTL263rnaxWIiVEU9LEeg5EBRH0d8XXUhOblUwf4Wr
JL2SmwkOa3ZopU2paLCmIzv2HulSz+FmDnIp89iFoyUhRwZVjKHQX3aNw3lIGy+7
9N7EfF1+woE+ph6j5DMDYGjRUoTFjqhn3EGuv5bv9RvirpQ1lQQZXKBnQqKp70Bw
EK905JO/gVGe004nibcjU/XmcSMFNTpNlVytcUMUpIfQiIzlOKj3eBYTOlEZSsGA
GgOUaj3KO+TzDVrFOwvkwGQ3T9YCuCEYs0tj/o43E3C4F4aRKB4ZTKRY58RV6Lh+
uFodSFI5KT05d70yEHnB2dr8xl5qGA1La6Lja7j16cV5y85kVAmpKn/twDUXaj3d
wXfnQngSxiPk6AfXMQAT0UPovU28a+bVNpBoYiXiGcDznXGiqG0PsRU6GdF11ScA
wILPO2o3LdCMwLI3aMJHxgRVQ8j+j9NuzjQFfjk3WiMO7gWE735aTxxbTQlsDF7X
b6NL98zfdlQq01yDynwD5xvHvaUcGeVenRaRnqxr36+ItrvmEzVjU3VFOBkDFrXb
fXZaLDefPOrvkJcOoJlEi/6K8CxS1oi3rQftJiN8oYb6lNdfXS97W0LGAeHwS1M9
`pragma protect end_protected
