// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:31 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
omeX1fkJFpupYOYyp110ose8za9ZBZ5ymOOgzsqHf1oRfOQ77STt/mkIVd9SIaET
a1dzOupkw7fR3QgzyphBaxYLlh0j+EjDDRKp2f/VD3PAarvZDk7Rwew5tmfc/KaH
QWl3S7u+SVhBW1QSRrhtkhRVWLZtI3kFB0imBkPiVWA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21296)
LZabUcSC6v1JMUW6Ge5j8DJJ1UXfm/5tIOaZap5/NNkU4QQ8m2lcD9jSa+iLpXW6
DP0Bamb6PyU6Ta24ak1p9SsOyNSJUtTGqu6ROZlv/w9G+KpVTQVIorqvD0/zJBW0
TvB4xv2IewnL2bdmIeid5vm9jDjCT6mmo4sgj8VfqiysI9An7xJzk+nm9s8ItrPy
tzCcA9Lz53btuL+AnGGpo4qTCK1Zwex+48rQLsrmR1NqSAMGaPYo4v4EdqfEvP+q
91IspbnXNaDdFFG+yD+K3y9AZHMbi3Jz0+oLA5GvdJ311MmZ1mgL2pUtC0dzpFKu
aUV6p9cRkAAwtZYMLcWwl6mD6KXxKuh7lZJAzUoEdbJ2G7o1WG4IjEVvLIG0ho8l
MFZn0/3NLf8TqFFsva46Q5cVQrcwJwcPM8Fwuk1ljO3kezH1xCYxA9y9yukx7FOd
rL/NMMjfNNYj7dwVemORDXCigmPv52T7tf9zBhRZlDdZEWQrGRAuLWiGAmOViM6K
lAmUWRqxa/jmFxBrG9mTqQU528Ut3nD0VUkHkr9ttLfs+jcX98CDcF0L9L5PWPJP
LgeC8sIw7mhbpZnalo55d5m9cAUzmU0MH3Ryka65KatzqqDp0QoKNXfxJRmmiSsU
X40HWFHzXjvIc3xCmVaX0sKKjSPMCdyl8mRpTPZl+LfvpmvHOyN/lmwRJkiCrDpE
YRlE0SsnrAEuNVzGul9LAHNk9BK/NGG5rIKEugPdlicf2Tx5pMXzfdcKTXYA7VgQ
AQbruD/zVhMGOpQ1bNyNSYZbH7m+6cIkmFlWxe+JFxGxqeQ1g2mEoa57oeOrp2Cn
o107l3rMhNPxDr/usqXg9R/lQEVWTrJLkhdhT/ntPcAS5THKbsFQm8N9SdVA6V1S
6q2K+F7OprPGN1avPLd2Kjw0tV8LhSYGwo1WQm2st4kwOdN7mvolPhTs204GmqH9
HGv8qPuji5iHOlW+a5TBDuMFg5/uetRllSXkpa/8uzbfJZqKINDkJx2EzfS58+Nq
sQSkknQIgJto7g9obOizmuAVQZSxfZt9XXGCItfm+Ue7AZxflS3G/abjBcARZrkh
Ij6k69xmJwdd5QQIyliVz4BVu/Fj5SaqFxqKInVTxQQ3hFyMWFyokzv8U3I0agyO
IRoW8Kq9OGhA8h1Pj70aV4XTKPK1FaFvfW5I0i2TIokX7tcUXrnEnsMR0lrSWVZo
fOkp04XvoAkV+EF8cfQsES1HjWzQHPvEAupvqrpO70MH+nbJ+boKApGZXcO2caIM
2hXoiR3nhINIaqs63YemUwyOU7QWB93Mxhsvz5xC/xBTTdXqVGlvnzAIq2UuPX/Z
Q0NDbr6QXx3tFhJ4vq8UAV2dqvdCozD2LLLvfSKRyNRbKo2YvviNKXoQ4k5BOFj3
7Yljelnxy5laC//DIiHYkjAJSXJZ3mjkNsz4Zt39D9knGbtHfZHYWeMCd9S8km8r
myXQ3ApY0SL4obeiu77JnH+viDJLcWbw2ZxiJLO/q892kiBgfTWzQVTcIfvnHJNZ
h6Rp9voOTVEbGCyDMLvvKMYjWgLf5u3yxYeUq4r+JbrMySlksIxITiXF+NSPZKT5
bAinxktDFcUkc+KpzbkM44SIp5Gft0alczUAsGgJhGZpdUFKtF/wpNegqSoMlAhi
+WwD681qWBnV5yQoJeUYNMB5SUJBWKyiCx+5t7t1gMcM+rebps23CfaqAg2Hji2j
ARA7kqPVWAZOGoxbwpOMraw0Sw972arwarXb/nipYr5jaqP0zYAb/3Ee4ZMh+tGw
OCESyRtLy0VWUSXZXDnoXqkSJhYyVuQvMbxNd+B5NKcAqcL4usO7FDEJp4ihBr9p
4dUAMryp0XptxwudDVscbs1D2LBFTI4Mx17idDXGz0IjeGU/6pIjViljFuK8l3q7
B7UobCVh664PxKCQPdiU6F4E8Amj4RsfFHdggmORajqRddsT2phvDCsHUv8cUeuT
VhDnexHAdG1BpUCzWGm8CyEsanRHKqWw2mPLX4JUXz68X1WgEsEAbIYy2nAd0bpm
FBabim3BuqHVGVsHN7P1HZMJe7gtvKNcyz4wuGwRowYOu7t1rQYWVPsGYKvOIBgK
4/OzhYnSKWYpASdfDUGHg9F7Q0O5JvL77RNH0X0PbAgcnlvcymOqmabDEW6T5li7
lAmcMya1Mcnx3YlUbapMNh1RAm2QpheoCi7ivmyxQZ7A85Fe8Ra3wx57pfIfk2Ys
P89CINZOwUMFA8vCuSRJHTcW6OIcWEDYQU7g823WxsaPP+1mWZ9FO4ZEEJcNn1JE
7zDqPSlgHtKaeS43HcSnHRiVfuvYPFElgc8x12Eb++sOwLbGy6FPzyhxNk8R2KOZ
Cb3I6NtziNYISyiBAFSI9dEaGXMjNfFlnukK2kCdcHbh9TZazvBP/HXCqH7VdLLJ
j4FE2lN3cV2R8m5T+CVJmyn/AsJFJlnnQSSfkGy0WbOu7WMWW7qfSagSjtLOmu4q
uEyt+JrgwgsB4h6ziLUGg0YpBBVZTJLDBhkp3TWtr59zBYeFSRzDicfck5peBVVp
napXE0DcXMwBmJUTUx0jN8FLriVXqLm321pyZ/re1SQ3tqajSc8ZAsf6WdyJmGnZ
C50kBu0zvx3j/ljjIVJmAF+Ch7hrI3VowHUUlnMccNUmmylv0vvLuVUJ/Ha/iTwo
pp5XFc9tSVu+iFHRnPGrkHxMLM87T0a0ULw+m0H+RefP+XA/4Db7t34GSbRpnksI
MbPCFuwDz2si81bi62f6rXy0h4v2vbnwb7GnqxB6wBbmYfZa3lRHHpgZCwhjVdiB
m2PVisGmWR3gUVX7vXuw78Lg2iFOC+sHQhVzI36TWUvG/PWUaFzTHW98rdZNDOdb
Sz1g+ts+YHJ9SQFykIfixlICBreHNS93CCVZN0gVKWG3xDzRqAZKBVyZ8q2O3bpP
+WebfGGYBBANDm25W1ZJjz79eFL/Q+JuzgqfifCwQ1RUoPpHSAQ2zyJa5uHGwCmc
LmSz34RvlFRoZxiPUmKNwjWiX3GC0seAmBxePUoJjC37Cf4JwgNkyGkFKoBAVY0+
6fDJr9fASGR3CU3AaE6m94hpx8ZlFqPKw0oFbtvECPXa6mhTZ9Zvjz+OGJBICrbu
gHQuO9XrOTy0A6nn3GiDWQZ5pjhMrtUDIS2bh6xGjl+e8CmVIp08V610LRLdqQWC
GnVA0AkyUT9PuvVOZgSyi9+1EsCQejaxA8UYHZoJPOC+XylOfjObx5OIyr1EcSJe
6SQ7Fk5vC405UMY+82mwMNnqzLvdWXiGuxJrixvdugqO5J2xAaH+wTIqIHsot/VF
DHQt/4cV+X+HJElCFQ3v3wiireZgVc0gTsn4QObjC7NxWg+QvPp42BA1u3bUDdII
z7R33w+X5YkOIyxyWAQ6ILtQtXDC1q2lo0xmLG8EY4xxrQqx2VDU4RWKefup+rtO
M9ckNF7KBy9ASMxb59sl7eXjbgCeNZhWyLi2L3Xi8uqkK3hsD2puCEd4uBFOCau0
RvUBeOm1BBF8P+e9UovrfbFafViEwPHqmvGmkmYb5sfOmyKhcSlvbxEpT0KNb9ek
LkOC/tdTGGOBYSmD3EWQLOSDqBgHSMgiMfIp5GrpYk0rW2MeJkE5/DsTpchSrVL2
DJikJn6EdG8+bn0jHIiCoc6XfshGmgIJpX1RDwp9Ti7vIJlUTaCz8JRHVeJUcHXh
NXp2bSQ7UcOPOLqOBCFJ3AHXLtBNPS/3mP2QvypUoamjP4Qfe2vvWuI4Oe6o7l28
3fdNa2HN+i6qjoIUY0N1Bqiig5DPa75LDqEwAk3TNepmPjR4E8+08TfdS/nfXf4p
buar2/etVgAWR/IeVOR6+J1f34oHEGfV78x7UiONAbaM7VcpJakGvM+rZZvuBuu/
wL993+5+SlDo0B8EjycLSiuGk+i9gZZntQJGFTVUSKpMPuKe4/XUp2WfBLEAoq+I
PtNviv9UKsrJDdgJ0xsLrX1tD0sv2pn6iq7lC/gYSA18xH6rLCeWEUraBcgn7DHg
cAqOTTHPfYx5jxVFn8zWoEw7kzRl6ykVokvGKLdSP71WukES3FbAiPNz/SFbseJL
5nyCrc3+CZ2kIYvkSLCfHwLLNPcqWSd9KnCXzvT82gM9kxNNZA0NsPZoSn3wQ2Uo
5LxJilF3t4vSlSDWOB0XSHypwOpbibjNU2/uqtRGtSnVWl48WYDIL7MkMRqWaTqm
872mba4Y0VwlKwFdi6vwzh3ZGNnGdASVY+3shkU82E60YPD2vxA/UEUJrD/Nr0RH
qL0csI1iXmr+vFft7Mj4PQ9HsxAWgaUIR7jQKlHlul6KhQGrelxNdiwX/gIwkk1s
T8uyOsGrdfoQnxrJHVKEPWZeh9AtYTOgRvYu5nyt33Kr+uWQs0F1KT1IOArkoxWB
HHta5F9FLAvW/N2Cv+5NqifbT0/82m/mlEW4NdFaZ6l1/W7eP0hnA+W8qvwvNcUT
KBzp25AQRr2nAYMDGUJ9r5K6yqWk7sy+PWj8bAcEXzZWKvfVaF77oXQar+2/ZVSC
KYSRZE7cio9O2a9rPOoeMSdP4eeyeJVvJ0O9KC5hqg0f7zI91zmsUAJ3nvpFCM3y
+mjbuHksRatXh4IoIUV3JaMbKyBz7OxwODhyJj7Yt0Dgk8N1ZvTT+l3Bx4cHvB61
1sF88SY3x+44YasRmERMcK3AR9RMhkYKa+Zle1sOimGToSRVBB15H1JW5x4tJ8d3
tsv4yeLBAVH8md2w7nKHIR/Who75M0CvYAIGEcRoi5aSJiGY/3NvZbcpSBq5lh+8
mGQnla4jS+Y/YM3iU4Pmej6QOasK4uKdeBy7GQScN0GdTQaD1WYwTSFqYmcqomCa
jlRLImOTA25C8D4sP/n4M5HoFFTweeqKdyK2KgcB4LlKQ+abovC0mLLCkioYGDVD
G72j+4BMNCqRUc5PFrjRB18g+3OVXtrrdmvfcQM/DkCOsXmLl7LWONQCllXlv1eF
dOkMJEpM2jqh16T7BfkOIud+sc8gJ/8l7wdkVKSZMqhaATGlrmLdGloeEwNAn75+
3TdgSzp0x+nNXAGlcCLrfjyiNkAcodDVcc1oiERLtGmy+gO+nEyfbfWIgSTO0GtK
fEIIzzq05SJMjHJR5p57zhm+Tmy65RJYJP5Vdx/VyPsoLtqJqwyWrPCeFbVJDSi/
fLYZP4Vb5WEY0fe/QKR+demRRCJZhmspiP+odhYI0B+M8YMe6q1Ux0shfz/qRls8
N2LBkc2o3jk+sVc7+ZTMCA2/zhBjlXhHvAm/9OTWQO7gmA2DwSeleuol4dtdOT9P
L9InqCOsMBT+BSUa2sGdJwV8dD9bBNfyZhMockkHyAODKOnyKhHt8J0Pub9iUZC3
x3Bf0EOg6Dd3kAAqdQ45IJtZNja4w7HbLZ/Z19QYHob4jEhCiISBBrZ9n1Zhe5YY
lKgufmHdDDOQ7KiCBWCi+2PCWzpldSDNHas+f6ZFVEjJD0JFWXw1GNNLSLrcmTBe
ANQ4NvQeARC7f+gj00shmhBKGzsflQnAwhx+QCczksWvTaBbKX+i6infCKRehp4q
rhxE1RrNA65uhw9kOAyKHlard1JZi8P2Assj0JWx6DPJyBEK97rvZDiwo3FMtqtD
VLcPUvedv5IIguP5Uq6oGj9JxqQ+8kk1NqDvyW7jsAp3OSKHS8r3XzMoDXGBLci3
9VXSS6pHzfmEYgWAqbqjK2rJ7NTTLWKSRk72keQiy4qD+Nb4xS9SW1tF5K+v/KVN
edNJTBaZ/cfFbHqLsebotC215O0bng7XRlOwsxDfXNzN+GqygBNIU+ymPEu81PWO
trUgWeZE26kmULFs9pfBSR8Od/yBH7xQqb4Z3cdk59YG+5LdhuTkTPI2XuFBIEeG
+jKibC3jzEQTIbduziFX9rAiSgotOVa5THYOBeewiSbZpzRcX7Ett1Stn20WiHeb
X6XliLttqzTmNbtVc4+z7+BqZk+lXJSBXRpWgL09MIN3FSqYuB8MsKx6qyaYHDLL
KgVlEz8va0R8yxniFCKEOSi9XHEjOs4Fjbw49h0HVq7ngnIWj7++EkJld+hSD0Hc
Gs33OwvzG2hnRbBKCDdMh+gSLb+V+nLNv3Ywc0WEVMxpUk/tJUi/u/+ozdmB5Ycr
pNHE+GKF15RQjQsJm2hZEaAeB5y4Q1HSKHWZotJDmFeERR/tJLKA31qN09RckOmY
SlgHRSKVKyewFEgFLn2A8xGNmD3+DZ2GtWbf0Tn0YbbcTGIcdAfam8tFOjBCm/ZM
RGFvAUd7UpA5cX22QPqWkFgf1qH+uPsFBFsAs5b8h58h+pds9jP6jnko688uUk/s
vWqkpiMRktxAiGABwdSu6luLEZLs8AI+IsxG/nEslma0D/Q79UfbUiKygqLhhOQ9
2hE8Vz3YHIno01gFGoIbQkCCMQhqSX1bH16kuCs68DB7T+7gymdDaT4/Q76ffOvK
XtWY55sBouOnH8ztzhRJ40Cpk9RaME/BHk6lM/U+5Ar/SOwqzL0762vj1/1gB5Z5
rxe9JboB13XGsmO9cktf57QlA/+zFDzpgn03iqVqNj6MfUgCJzODZClYukx46afM
5A+/BvRS+3611E03U4HA4U8LcjjzYIpHIXN+QKxWs1HLQLpxT5C6HusC5h9jV42E
Sae/H/pB0dp2j+5ggCubz3aEjbUqZriL/BDaZWnJ6hLTDsCFOwHNP2F5JL+dRAyF
W0j2xsZqSjkkUTbActwYiytduM5cZgFDMHRIESAIljw3vX8bWzYnHzeuEzVEXkDZ
NuFmC1zNOdNzD0jMCcKDmTZGaFGDzrxI/m5R5+NsQL4lg6WD0lS04og4Xh50VPah
B3lIiBOsAGRQsmlFAvDSPu6NuHBa/GU55nEbhHCpNSt665CPg558m3wkc18eTHzY
AOIb0VgcxQSb4p7YgHRblebaht1xowArhPnpP/ZxgwLlHA33ZmPEeMKK4kMxsUMj
MWTRrMMGM8lXGDeYSEq8GunFzUQNdij0G/h7fSNGBxRjgTEwGKlqzvaovz3HExFf
QWC4SF4/Mm5z6eYVn00D99WYR5vWDYBVmdwOoUzju0WrQBkkAbl7Ul69PzdIm/9B
y/xUQMAouup9rKvqeyHfYGCto2n9sQY0an4njIzxF5jdBMD/vNHMJ9LvscsUzC67
zuS5SUVkB+ar+WKiPEhX4QbWKYYoG9eTPYMJpw2iu05HKT/iPasMnfgzjwTHePWp
5rJrmmgFWCvcgL+r2NOZSBOcJRpg8uvKOwFUnZ2SPimS+hJ7rlcQhAza7UmOzP1O
26ZUjKfo560+YAWINt6C6aFHj3esGU7Yl6plkFeAk2d8Xv+hIByQirl7LNQWfOoQ
rspsNa6SskCgYyaZPEx84KvYR1Mun6XN4g/JsbnXI3nO5bttLdWKh5X+AMjkFkBE
YlCX2/Up23Kif8Tx62QQYqFaFQ50bU9Ofa9FaGvaKtUsS7auuuN9gexpgaKUSDZI
GRHSPnrzOi9mswRhmbbrTU5nHAZ1BelWtmmvbqfJCcD2wvBX05Gn75LgHpgFh9pv
RQnqmiAXrRE+dGa3GNSm8e8T482Icw832vOnP/i1KJf24+c/Tkpcc8bGTUziMFbI
oqc+3/D3cmizx/rXtnajun/AwDekUBzRN63KEWSngWY/X9k0IpsHh/CL7o9ZoMxo
w5t2svkDx/s2LfZOLV4AEYPeFWkJG55Pf0/B79mfEt38i8Pi3GQPjCPyax8XPRb4
+TOOrL11+Bwiqq/26JdMVFluAFLc4Tmo42u8M1j8MvopPTIoVIIyT0TeLK2xtUwN
wgPkzInn+2dTQ+/HGpoB794lxfPyxFqHN9ayrZ0x9cDKSay0fTF0wfPnpMk+Sq0e
jKgbH2X8nT63e64KSyovYW+6pIeAr5DDMHFlBLUFQ8pId8DjsdgbXLkpVvCZ/60n
7Shh2lyC7PfDSDqLrsD5l5XzeU6yu6CT7qFYrrDX2pHnswpttEQdvnNjTyagFLm3
a/Jo6nlNr8qtqRYFauj19pfkWhuzWLybfvRVwQJhREGgBbAq3WuRj4YjxNBOj3Vj
wm501gyugKu75QQZF7hGb893m7ZC+ffmMZQx8Vjb04tlyZkXUCt9JMf/hAtJsrPt
B7aLZG743jijTEj+nKPOn7yf/BL/AXCrHg73mNjjrq4+zbynssUBeh/spF4FgbRn
GRYz/MEH4Cz8nJ7iXw+DKTPU7Jqwo50M/UDJp7x72egJ5AAyoZ1Ef87jk4K7dBjj
sUFnaZXHc4n5/9lkF4n8WL/uYSLKKZHrVDY5zYsnHwB7zHMmXnRotiaVHYxk611u
I9BFpTtLdA+0BPtwmbnqVYJOmzKM8CgkWFV1KweHhmPvjpkI9cGOHie8HXLupP4u
q4199vI/bvRg07dKDIY6aDvOiro1D6nl/vwiDfiIFms2zHYl9XhP+aRK7t/LPQQV
kLIX/i3iP6aJXp6E00nnO9sJeIEOiLiRw6yZ07hHV200oDqVzKtjsSVzm5ndNHrJ
QB6xE3n04cSJotb7yR6aNa+rh5BYcRO9gvfZQFvqaec1ESpab6i8AnTf3SKBzg3b
oukQ7K5zQ0cIrXTBXul4Vx5mbCUp2qCGb/7MfoIwTm8k65eOEotG4tpiPIxVsmvo
3zlMdNOPmkWQGVUy4kVE1eWTQxuay1i4TimtTKbrtY/2cDEZwWRo69OpmdRsM0xI
qFAG48h4XdNAH3iBlk8MfWtBLeVkePu1QJ2iJbkbwPOIKx8+IquBq5v8sQmEeg6Y
iioBerdxa4rSmhhK11dXKFlCr7YMLwGtE6yVJSIFvTx2gxkvoP9264cIlkPjuMMa
+21U0ne2p1u/BDOoT95EcGM6kBhWNsS7Q/AmwMwPMwpzHQyLTwRaXWyZC3fmZMUI
m71qlHJMcUvtvCioqBn24uZZAt0rNKSNE3zYO5hhmcCaKGAeUxHHipCRNB+rvM4y
ReH1g966ZzzfJhjQFQqrgS0yRq0CB2CtmRSoUMqB0iYCvnVWEb9L8FdkKvUf/Czu
rYdpPe5jaaTWkaMUtY/zrWw3Zc8Av1y6PIVV1l5k64SVr8XB77doit2elRMRRMXC
zrQ/+Oe3n9t37SwRgAzGyEUB8uxeD0+SadTzCU3EtZzZhtE47EZnWR3O2eDmv4Vb
5Jlw/JBIJFd6dwdpxaVjoXA2+13lcPL38zDPakbiM4zcc2GZp4Qx34gkWdhT30TQ
EFv9sU276KU3FNDEC6UWLnP+a/lsyuPHGhfYoOzd0QvrJvbK0KoqXHf3yvTN3WUX
Ywv4Mh/c/DZbmIbf12C98gaIYOHL4+y3QgDdGkwQWWoD8+UG666eU5SAun8tXxTY
7TCI2IiY1D++lvFpBJrF2tN3cfjHy/oEAvw5NpWsLXM9xDDcHTWf28Olgs7oCy+Y
TigCxQqZ4Hl6XUX6BzRmYYTRByepivd1P2CNrt5fiwtXRKqO1zFjx9e3Uy5jDncX
KMZmNhEwFuvvQFT2If+qlHqXOvZC4hItSgnKGikEyqMzyhtQC4SRJe6XsSDKrQ9y
hxL4GdI1VR79WVWvl2p4mq+J2Qm90skO2zddFZ+Mlt8AR36tfH4VMySQwVW4Z+k2
iYT8bThyG8RdD4UvtSWSRO/7vW8yRTjeCSj6LD6LjM816jbjq4UulGqxDRvKxFa0
rjm1cb8h4XARCe0l2NnzBwN2GK6IRDAWlaGmOqbPWbn32cqyrQGqlGS4qqzb67Y1
2KaelssXAKebrOb+6LM9Hn4Quy7AkgUn/sC1X7qAc+r5hKFMVjxjcu68LoqHS8eO
Eb2QgBotK1Vkd/AE81PM1oINoDtuW/LpVgYOEVePa2Ee/UDaBpBd5zpWxaSa37Ug
V9YPEupbzZNuLGewNG9MM2OnHlRCwPTT4hM7OwVcx6WaFPobE30NSCEPNCrdwAcB
1kkrBawzTGgPez66nPgQNdgYNVmaABDfo6DAn8JCAadKNCaX95u31lWADlKo7CHU
o12CR/iS24YXRyhv1c+Jes4db7aCUPE8bm4hskNNX02YLSyee4ION6j4f/AMuu7Q
CXzVlAbkUF08WXgbC1jtdOCIUcpOGgzQDlOm6CMYRGEoDDNi2g0PNmxG6Kuwr10c
JlM03j/I/8gUx2XA6qAC1ZekwwFvAE9JZoKyoSEm0QpdbYeq8nkolbr5fHaMSRN3
8mDRr3d1LMB2oGJkT0JK+hACyRksDnGKQb1F2uGcgErHqq8rLsXMRydROG2R1vyJ
5+4J/NcuUjqXlpjyrZImA9WBUbsG9w8jZgt7Ej/bUQGwJn6kjms8385pSIumpvFm
HEOjIlK5SiaabdPHGNjLIj3g+p71NS0PVxn/QXiIOMz3yTyRVwPTy7WX0ND8lWNc
8tVSChszzC0AqoQdg8nI9YZ/Vx54X9nHjW9zdd5xh3IDacLJXI8hWtyF1xHxeHhY
2IjUaJgQ3JlFmNaCQSNBfRG83iBLg3ZOP4rf+ooI/z1dZGMsdiILmlRfZGR2RXJW
IV7/H66RUWxdZ1xmbAL+4hI8gbFsd+jo+g3LcOzZlb/vs5z2geWeoN74h0V+LDJv
DpaOFg89zmcbT5WUlXoIzvGwaCf/j4rZienfnt4pk3qr2UAkm++OrQ25loVv0UK1
Ud+HHtR0DMMvGEk4eaAeGDXSKJbHrAaoVp7XukjnEbZsBWiuittIkUNF9cZNLyPV
eM7CKotq9zGJlZTvs6bWI8a7a35HKLj4kFDSQ1zIOcvjxGfonbHBjVRhNQ7g1ybV
+e7FPvoyOQ3Sf63o8mQJAh1Dl41AS4gUDspK+auFd4nC/DbzZYPDi6wkpZLpuRu3
4j39TSc3covZu1JPDZuW6ss+7k8wqehqLe4Gafxr/MhYINCbCch7bXErsUjZO0DL
fVYlI0YSC/PRwmqWKk0aMhFQsaoXUoWZgtQtCoLjh7fKI0RL9+pZrgT/NLBshizG
pSmE5n9wxbJoL2I6l5CZvAn+yc8jfs46T/WRQ/6ZzxkD7/XqpIAoCVV5sQoKt9ye
5iFsWXLPNLyDgixNgCa97bRSRFCAheazhgkZaR5AZ3VZrywsPQjjC1YeMCK1kooB
sbJ751RQ8f9EoHZKGhHVVWXZ2JHeZc49Ap8kuv2bYIpxHstZQ2kevZTlWvcHnp+U
WWLhwIdFzAyLKxgj5gGT6fntGR0D0UNsdmOAdNUUppc1N2s9JUrJYsGbs2Y8Wda+
n/f2pGCRuWugyf87hJX+lF6BU/kHKrPD/5zPOHn1vk7EGVQ9hD6pgJrT4JDhsQzP
MTgYmTn8IFMwZrh3Tu/k76vMadY+B8mj9VEUvtT2Lu96zUYy9wQAgw1Jh7TQI4p+
g92PLmc9IsdeFcpqnSwCyKEEnPaojrPLmGAJ/g8xkXfZ7LH02FjPsZoOPKZSAk+m
H4zhRbPWAry+A3zMf3CsHy8i2yvAzqciSI17s9GxQUNuMtOCiyCHl/BVhfGYKqy/
oETID9RRtNy2/5V6ndv+z4oGeBEOkl1Oy+doqn+kK6OEd2lWi5G5xoVKrbCfnhKD
IHhb7nTH+u54XMfM4zE6CKamAt0KfqKNAeqIkgZa8ag437KrwuP2Twc+d9wYYSm2
ElSiIZPFgBksbDoGTsR0R+5GG2je0K+xJM39c9JtTduFaLHmVTKkIyL7SgSVBRPB
+IlXmNa/AMiCM7hLNCluHUsc3UnoMeOJTMdvqZiqLCCwruHDHWjH42/1nk5btdf6
fUvuVBD0sPoQZuEzSA2CRzmYh8WDnvTbQkF463lPqkmNKfg/qE5cC/SLqQ6p99UM
9y/Vms50vw8JDuXU7rhbdWOvBKvDBq+zIpMOt5RmOgQbGLIMV2Puimx1PWBKNy9w
PWuwJrPoINXOwYyu921eZKg01zZu9LMkYjYuEZMfN66Wps7u5D9oZ7ojeUj9bGxB
Icnr6aTHKhscd3AMTl9c70t385qz+BpPgvfRUdS8c6koaX0YLZe5pa2iWMWIAxaa
aVrbGIbmlSbXGQVTUjSdBvYYWrVcqiWNfvVfWKdz8C9OIPIFybkL/6V2/L5V9ksz
W3kw6Q6Q0WR7Z7b/QY/O0jUSadF7JAPVVaVqF+aiwx0Ug5AHqqfgBohogFXxTNK6
ZEl/aM2GavEDoQfYOjsyzP74ciaPjot5xC7/o/0uTuACuBPkfk3O3HYPIisgA9de
zQU7neTU0PwjOE9X8lAhfGMmbI9wKa2YoUFu0oh0mSilw+/FeVr5umuijNB+swTv
2ntu0Dbz62wg4CGUTKheQ6yEltvbK2NhlfTbfbl/VO+Yahc7LbFNc8fYFnljZQi3
ZNC3r5hWgmqcfz5GJ4S+6OTv5ldg+zc0WVEPuKoeX9JkcnzvD8yeRT3x3v+vyr2h
8fQ3Um0upIiOufuc2pgf67s0/sia6gOrVvDPvdpU2HbPItdg5MFH0uFMjeFniJBy
zkgQWFNRnKf7F0sREmTsZGObkQ5v9T4vtSH3ekjVVPrm5IioEe/L8uoIrmRaOH4b
M551zNF3boR6XJ0hkMnlV72YMdvlJKOHgPdGZT+uLbCcJ9MKYBFn+/cGDNlkVHku
pEhAysEpzD8MmYgnctKEeWKjlQMQKchQrw0TBDjAb0oCU5K8QI/cWaBgkPmx8wIk
EjxVRrLpmE4RbgMx77Sz96ABbVtrDqMLct03mcdqPoogzfgR8DzVeUazj4GiCNC/
6ARp9fITpHMBmv5PnWN+CGpcnE1z7gH0cOM/uVQ+AKbh63Ky51v5J2Bk+hw4WY6g
QCjGVVrrBpvCjweApyT8hMrDQZDUYHNeW6WMHeS97edCP8IYUT80ImuSc5SQ9y7D
SQ8rcAxwlU4z9KwVlnaF3d8KpAXv0Y1WzHiGsTCnoj0/Hbcd1H28m86V6zKD/ICe
sUDtwUdNGHQI54dj4ZtmEp6GH29eOgrhaMjg2ey/DMrKY/2hIuSNsa/CO0gnflaE
XF/4lBUHmxGBR8mkRWOzlqM+fr8QnaPbPANVJshRsxacbHwYJcjT9tgr0rRYDWG8
0QuOI6He0x0bRS5r5jR4cGlnLSQW6qMeTrBf3qjYOHuFKTr94zYuNa2s3hDGyhDo
6uraaRavgQL2v+wCkg0uqVaFcniUixiHI9kViDLXa8O0yk7eq7RqDkmIwbHPZfg+
Zot62Q1plT/+LP77GxyxjGg546CNA+Pgepv34Da7tFULKBoZa/hF4l44glJh7Zqt
9Dyk4SPhw4F9/0ru241WiC3x/agw2vzs26TVnVfhdN+3H36EcVBw3osy5iF/Chl2
lPuMOfytjjqxlGFHtKlCRi4pr6CCAIymiHt/uXtAJDYk//KNN+xy4LgRaL8466k7
imfYDMPIS26eprexeXvsZkf3+6w+Zze9yGUjKxtdbGCLg/Xx2PKjfV3Yi+B3fghn
Ti3g9ZYRiUn2UDY4YE0rZEugswEgcLyu8PgSjKzlVmCTLCgMsQJdNIZ0BPoMXA8n
9gVA6Hi2CLpmjibXra1GJNgorVazaW472sdrsB6nEnMNt+Dop/bon2mKkmPJSmMB
3GDTBf7FyE+7qWnzWt2Ohph5N3VFMzzJ/PuxCFc5r2ccEO6HrfY9QLV9TcYeASES
QXrSnjnaHZHRoIU2Fp8e9NZEXK0YXJgWjEXux5PPyVHidwr2vZlUUD7xo/suPuH8
UddzDiFkhhNw0BGOfUfi6EB2alhtTXjoMY8K8jVPBb59e29hnumbgR6bPL/2EfK7
ZXX8JTX868fw6j4KdwEz1diUdTMF6WoUYlAkz/HR/dcns5AQf35P1r64ljHrcb9k
soy01Yi0epFV+SP43ElzDckPFNSWxwyWNBZ3P8TkjVjs1O0LKMoIjzRtLj5/FPTV
iMkuxx2IqFInewM2SQzKc/xa/FqEUdrNY2Tgn+QKvKOZqV+6+9kXDWAvfvGk2MyH
w0uWUess8ez0hNgzbcIxT+DEVajWmXiI9V6l9+kT+lC87hJD+b0HUeSoByt28zgv
pXrsHM+51FvJQiqsceP2H+iLVGzKZJqHXosxJfbEdRDHmmZR4+uiImOaQ+QKSCVm
vsxcFIWOfiztyYeJRwvGCA7+Q6avHYBZ4EhqcEdnMLuz9Sw+FUDAOdB0GyJKRZS/
o7Jpv05VqdOGoO2rEwo+E2Wm+z+84aHtksickp9x1TDEX97dPk8wcCNZlCfE0iB4
6PvsMEzk51UeXK8zih/yuV7i8fwmJK64shZBrd7+iac+3Gg0TsqfVCSU4x1nmhru
CadQk50Ha8K8Tcagr952PG7cUUJnnmrYcK6XL2sgvMxIzu/oR9BPDX4fiWnzafnW
ackCrFadKDambwoHJdH0S5G4pltdbtBBjMDl432O6QtYPX0iI1gcQthYGEIWukY/
u4E958K6Rbwcfb5rT14HUE5X3PFO69PJLF8cHhh7ZxM7cl3uPc1mXHE4cs89ZNGZ
YR5qh/X6qwr3HjpEI+4XMZzjoz4VRN8Y7XzRl+dwe+0DjqYH4TB6VP6sVOc++Trb
CCXlwqiap6ucBWVzFdaaklUk80RN+RT45/OzQKBUYZVZFr7kHASyGCnFSKH+dQB9
z+saob6i9wqx8jbCVglSrURpZhOjaJYgOGI4wAzrXqmZ3L5qUEc4lFHoaiM1GxeL
zGAiLUl6g9gQJB1n42OzKKew3XTkYUVDHdm1ao1sLLIqoyFIRh3PxXAELF8dePKQ
y6mPYtkUmjeTGPnYFSjP2svVy6xWyvWd0fa637+USpkurnnBdlc5mIny2yvceYjB
cJzRDFqxbOA6DxsKJjfL4P/AQkBUS7FXlX25SxEotjR36dq47XXz1lH5Y241CfVi
LiuPoM55SOm5MY80LoqgrO8v8slc3aqazyw59Nu5qimwEMhrFJRW5K2cy/xyXPsW
3fErOpOcgtT+Ls5kL4eHK1O/ssXm0ga+VrRKmFNgxNmfizqE+mdmwKgC//p7y+vS
/ycA6kP8OxL1wUWqo+lLraPvWMMCK4iQxWHWokNSFsn5Gj5x3/92hkNqclAUH04f
RDVB9UdgHa1UT0bHN3recch+rX2Q+0osx1eLwxJZQPX59K2g5VRWlW/xcly6hI+o
BygEQP3fmU1bPcomLI99e1Uyxautp3//5TEmiHZDeVmVTodRFEFK0Wnj21WUeJE5
zqhYEy2uVFTEVx2iGJNdUdhsofAVBUUFDcT3+LhBSAH38t3WWZmU8uwzF8oZNMU4
EEWqexTYVGklayLRYSzUHLX83dLvBYLHNF7xZ3VEMi/Ir0HnoIO5zA0oOQbGmtUV
SrmEQ8FfLa+Xbqq8ECC0obuGA+TpZqwgeG/KsQ4euXv4rOcKHZ4lyUfWn70BAmo2
MK1iCnfb4BT90/KxgoSsnvXSixYmDnA6CGN8PT/LY115AaJir0z3/TbeLI9GaHVi
oj0mIO8nbpW4Lfy01NAbsmPUKTc6yplbmpSfld1Sqr3izmdTIHuZOb+CmN+LQzQa
6nV0R/IYsM55FDu3jVydbQgEaCb/F2lWuKyHQOWKH7yDyz5Da/2NeYkcxIENa80k
kd+2q+Uh546QcSnuId7fm5uMFcni85NJi3F+70BhFCKDvhbdSzSi31pKPWBcTKpV
lEOZQ1ah02QBSCuLJrNKiP0Sms4abvylIiprp4MdAxxEHn7d9K3OuScPs45kwqwJ
EEICgSCW4gZZnOlfDvF5K7aTJVd1mQPgVc3t9hMZL7gF4z78zweVPCRqT66ib6pG
GuU4N81PoP1FbnipRVcA4ah++yfUG4giSDUO6ozJYwQ6SQrTlsT16mYmd5HhYSph
ddGOTRhnJ7lf+f8iL6H8fg1j/dA7eVBBOLz/PFiJ5sjemmw7avfEmNLcSiNBEOdK
QOXwqsOxr93rjJaRnB01ZmoXUw19zgXyCSbyDtJSR+S1qOmscVHXGjgxfnPKdncl
yXCDAgCkdU+JB3CehFcNDzVSS1hc0/XQzxM8Z8KaOUWbH72jvBSL/QPCK3xB2eC5
qQEQr1apyz00jg11HUowjLDiZyBUsyD4TcF6JSf0YMFaJYsty3HzeIdOShrF5gsu
O9pW+nRVWRHyg+wluQVv1b8gpZ9nX/ZbVwHFujKSSCRrjwqdrl8a/PWs5rvZtm1c
TmtCtLTwxqIsgieVqwDfUfzA9quhrpFRsZ1aGh5jirldEvwTOicSGqtv91pv8iFa
3WnJEaSE4co3L3sCFb3OYCJQecLjyXjzdxrWslBC30Sco74L27BLdCYx5TEUZsO5
iLl9YR8L8nQ5ReSiNpuNOZt7kk8Vka0aflGFbCY9rhC7t2fhN+nbuKp7rG3u9Zxj
iHx/HCDJoa+HyS2yxw/fFaTc7EzKOd5rz6zu0oaWmO0HPqvXPPBskjS8ygWNR/WR
YnVRSB7dVCjpeK/gu3W1rSGt7wmffU1PTpm2dXEAH/fg7lz9S6sUKWQhyEh6a+pK
sdYGV9cYqTHV5yfUIiB+1rFSjrdPzv+xiCzJWOVYPbkS7YE5nD3VfIQFbYCdOtwT
d5jBGMI9rhGYJc8daRJQHoUKJ3nKZzm/kwksa740h20SITM4Sympj00oqSmGSIqs
n1Oapl9M+JDQa1HljYRB4K+EKVCAs9vdoPDo8MBm9ZWJDv0kwiIcjz/iROCGLOOe
V4gCZmMrngGyu2LGrGBHQDVFDiSjV7PEi3FwgCJZyh/rbhIzywlmvPOvVGPawN2W
QY22eciC8MQq4tgXHxBHy1bgFwL/Up2nAKqC2PzZvTuHp6wW4yjx6W/RPBpwDHEO
n1nUPz7KdnIVymS1NsnkRoeQxYUQunIWuMCz5ZXBrI41CF0Qe8R85tMQZvJ1DMYc
F51zedFBuMudg0AYmkpIN6XugyBgYMh+IDqoCvfLh6QrREO3vRhwB6xgOcgMLOkN
6BqdQnQZbvL0FV+hE2zYCzqEgvCQmwwbX40u8D4CacU5UQlkBApStgg/04DgQs1u
tiqCDD7rbWjuDaOEEyIpYi6zWhx1rTx/XHlj6v6Kyqd1NvBBU/iyegNNSeatdKDw
D4Cij8OLfMpMgJF0HvyMxbx1WdboRrrX7FSMhvFIEORGeUo4z53BijuJuOB4nAwz
1F8tm+XnmTD3X09GZLa1W6OGHvVzARm3OTqzdc2HBVIQ02wmC0mfi/xufHgZcYWe
VjRT2MCD8ZReNJcabz6pvMLLRqZdVCJaQh3CeylG9/Jr74ePnz/btn6dtxXCUC4l
/mMih+T0YraEoe7AF04TnWmQuEu8Xas9GpOcEK9wYSHx+XQc0ZVTUidk7gw+F5GI
n/9pE8Hxfnkdem6RWOUtuEXaCrlQr0RIiRE3TBVDnXQ6d38J74fjNOagvHAV/uc6
og0B59clDICuRXAqKkQIit/Yf4fdvMTZP9Ke56kQVuVGiu3wAzLoK1GtvsLE8S6I
0aIYEEPiKUaYgbd5QWCKA1QqtJIyCDBtcsrRU0quCXqYck57ujN9f9+mdVdo5QWv
/NLsNtbWIXPjfKckvcZTNOcV7u45QUxoeZ5bxnOG7lJ7oHE5MTOX8/WnR7Ph82fL
ysK6xFT5hBanCSKe8DwPA3VERYotHGZDshtt9k7etNs4ZQROcKU4s0HP9v7h705o
Hag02In9pOiIrCdAIfKJsm+GVeWsDj0hE2UFSb/wyrIwmwwFVYgwTeQuLQUCGx7m
1CFeUEK0fIhuCSAZNmkmkp0RKZqAXZ+K/BMk7X+gOTthkj2CSK38Ag9yDytvRZeK
CqqJSYhF2YbRS0l0egzCamCj1ed3TZt0JGO3RDN7A0/80w5q45YxDHGum0lSvVDI
h3DwRjg1XdhM9D/AUj59hvQJK0GLZmkY1N7cCgMko6Bw0MMfJFJ5aB5fqXhTJehH
3tt2GmzqxAJ+SpZEFDZu5sy5xLFxH9ZrB+0IKdQi6lFWc14zWrtXh1o3/ccpsIaO
PoZYNE7Vh1IJQdHcd3h6uQSvG6tMU+xG3Bz/Sq8kdeVVq95OgFQXVVfAPdZokWOw
UZdH6nznYsLqxKZ+8DobyALCjvB+jqlHzCRELqaA09n6A8c4El8fDnuMU2VwZH+G
vS/8yDWIGXcP4204RYsHv3HQFkxYHe8gBDTJbnPctGTns0oEZ3lnTmelLll1nCbA
WAZs7rwVxpsMNhPngGHDOQ9/+aWjzEE3hA8e/vgjqSW+ugyo+0HQtEiLI57d4C38
lwo1Z7V0HNabBuiWYDKJeOk3KCBqpKAtQlTk1tJsm7vfpxhRCqW1JvwIs1/hq4QW
hrjnNrXc+q6we41aMIdrzYvpqeMSOMUcl2WkeDlSh5+mzMc+YpvEV9os/v9BjFW3
hcWYLnykkx7nfoyKs5mPw9VQTR66MsjNIPL49EBNEbew4tK/03Pmrcy4Gw3ZrXj6
XPdg53JFiNcsClJoOQEuaV8rfcKIYIJ6WGN+osHvjgthCcN2AsznY+LMiFJPR89k
5RNP7rg4jyqE07o52NJaedS4DEKevRD/SQz98RXzQVeZWNS3l4S31m4xzGd2GOsW
tseaC2E6S00pQd4j/B0oziDqGDfjPpQyXxE1g1kac6xczMweTZWMCOfvsbCGnhw9
npZNgUXLrZd2t5Ek04ihA9sy8WPDqQ+Mh4Gbykpe35kVFs/4PmFljtkIYvb2se55
E1pzWnwAB5oxvz0W/qFl6P/V7AnI+W+kpNMdbJfM7Gv9tZMyGsQh1P7ed/ujGdc5
J76ihRrg/RWoFmobmCs7FeVXR1pmnnLkN59c54qguQwSloresS/PRgDBX/4qY5ez
4psYIEEN2GFN6ABVEioXCL0bEw2UEFVmgWFTdAxOWqozrQd39SqxWaWb4p6g+1QI
Jr49Rt6r7+Wo1TCwMQhusbo8JK1JsUHthtrifJYiEDwKt4+fqBKuFP6jA2SiPrJ9
N59g6SwJTEuFwTtWEkB9lJxrhJVAS71Wv/zCw80e5ZtmHD39HbqEwDD3vAPCA0ky
uuasPEuqaJZQGAcAJ+itTSrybTsYofH7p3JJpYoVjRL6ZaBo5PnhLCFiczaDwTfJ
HcbW28y7EFujLURYuHeGMbMOn4sl30h842oiY3EAVrYnzyHxhWexIDIuROrLyKkQ
L8kamMELFLoOy85bxfPAvsjK2E+rTSa7411sNMxWVomNQyh3I5/Gg/mt4be6kvVt
WX2u2iJgMKXkFax4/KMBb4tJIFnDZXWBSQGRMO+QuC27LRznDUVUnfIS+dn7uT3k
97gBmr86DaaCARYFHNk7OlYUXWam/5cqMMbmSv31SZZj++md6orkBmflkJdDhow7
6yuRD3TqJTcrP3Yf2CAkxsqLunNRBYr65OyQQxhil1/gLcZWT6UZhJQaaPrwpVEO
4kwHJ9p91h5zfM88cWi5p7kn6sNYkdEDGOUGZOlxlr0FqH3AsB2oykyoKXxnPveC
EiA85oYzJzYC16j4okxrI/0pHkUrnGWGochgVPLEyXB+hHM6dU7sB3ZWi65ohuiS
0y108h9adFcwZFu14/LcEtkXQ2ZpZpw4OOxOTPJXq0fBeYCBx2AEWMPfdVJziO6q
nBAvfXeHL5TGl6CaKmo+7H6H5XMpLMgHHmeWnZHZp1DPnrb4uzM8Xityv766Q68G
grlPV2RaeOQWYZx+Wwac0D2xKcEVKW/txoGjnzjPTAjvU2IeWC0IupnjMyUFEOAY
RixuEOQ+zho6RSQWOcm/JrRswWj6kNJqPzpEq7IxjEbC9813+2Tiwx0kvFbOyQPA
u5EvWSWiNqJkRyOKCZI5uwtpFnxMIYmIuqgjxSF+yMIDeJC//6fDqhZhO28OTQzd
2AZoIBDlwXenvULKPgWiUJ2Q6WFOgL4NlQu3yJYbAjsQ7kImLcjBW0j5KJy4wb3q
53XIwaGMtw2qJydYt9E7dTvJpywsWUyr5l6CosoqMue8vvvfZFdNXGxokK+ZQAXw
gKuVQu5Me+pQMq/kbFHPddo8xYx9GfwtaUEow0WlpBqQRTAe5aw2AKEajsDO18Gy
hzwnwx53CGB0O20tSeluNnF+0udCjX9OjzPMx1EeCfJTG+Lo0l82WKVMWrUGv8nY
RFYgXoJtd7NT3Z+3yJ/IXr7qfW7aFtA3XB52vf/ZhDTNIUzQfKhocH9wwHyaQAvJ
OvjUpnW7SwIkeKhA7nNG4QArw0CNeEgH0yUC7t+Km9zbOvMqXsxPwH7OJPXEiHfb
tW/PSD6AueLg0z29gVa2b9UQAZZClaqha7IawFfykpEwowIGSRI6l0mrtGgNrJNy
+AKrT+bqyX/olbcFmTpSDEJPD04cOHU+O2bwLVUMrmLh46HM7Bw++/33RBnaCUZp
bK8Dd21tqzA7lR9WcgHWJZWCNct3hV3CuGvpZEuvYI9EYvnU+o5ZaGYbAmKM0CnS
H9HwdViGJb/V0k9R+pkKNgRAfHZosr0JLIscuXF4aSsMqr0r3lvcd+/PKsKWHI9W
Ajnoie7Q9EBWDeH+TessNsHA07fkm4A4LC1HcBaOf9zdLTSkTSRZNAtaL+v3QaWt
W0W0WXsguS/lKHSFN8fwX9NTi/yIrtZhOuJ1diZUtUTwxuZQJyy3PI3cwR8HIBfa
QP3haHaDx+39RFykeefQMYlDIiHDGJ9EFYe6mxkp7nEWQ4P6dytFGmmVmEeu+KnY
HjZo0lCcHLSqINVzNhPBLzL29R6t5QNlvCYJNOK0W481qQxwD/t1ktm8WClDXi9u
EPaL5e4zCGGdmMFY9CgcYF9z5kKp3YJ9lGt9H8AxbjjrVEJbvfrxLbQZ+fPSqZ15
QLyeG2x9ZoPZ0keTIrD/jedUg62tyWPgo8zIA/ZSxa6oJIaq+5gsl6foMn74po/H
Vq8QESRLdOuQVINS8M9z+msmN+7+qXEuSeKrOoTBYrS90ShtkM0tS/WzLna+/WkO
Z7eFy0tHYIEODh1gEsLmJVfeKh1ysZWx0sMl4/kNuzq5TGSBo5Ixy3R3XjRBkBIg
0hZ4xujgYrV5vl/lzuV3hbafbXITkRkEBueHMPCADPSN/ap73px0WHDmNqdaZWAA
oVhdc87GNQK8JqwGMZM5onl5ZZtGZ/4SXcGIfq2UGaJauoAXtsQK1oXAopwocHYG
3f9j3cYWpB4XaFtVZ/ujSgQD0gdzpWw4TdO7MKEDhpZpjHA17kxeZCguezD7BSWg
eS87itwL7CDswgMiaNzXE5vgK1A+7AbneyekG5WvDOXcI7FFuoApP+kNA522OM72
Bxx61pR/tI5Sl4s9uhayBprs+pRYY6GtbcudiFlXB/C0idIN1ybI4TQo61vfDgaZ
Tq4CeErRJV3ib22RRB3+FCzUp3lUKHjietxXe9E0+FUKqemQTXDl2NJXPxGjcEFd
kdpmPE7AnD1Jg/yyMaRachwTqk+b1UwFr7qaRCVH/cfmpjfPs0LeVTI0qGUYz5vT
e3mNQRP9BYyRBWQ2gHQksIx6s3bcsyUVZ+L94ahfvkBNWrCfUMoS06dI4Oy4uPMT
F16+TdEPMPbSA8PRV1r65yOTRLy/3iMt6AwsJvhUU3bg3ELahzZOcbfIn01XLY/L
W35DlHCVhjuNcxtTUUzXLnovtnz1FXTa6hj38T+yia1x5RS/dPk51vfhNT/v/jEJ
u3L4qy/cfnYsQE2N2OIBVwC/RmFxcpLrykFSJv86csi/uCyHiNEkNn+uiboGwohX
aQ0RxpNiyc/FKJOBQlpeEenJgpRIoB2GRS+T7XV6X8Slevkk9Nb/ELbWvXmjJzwn
bomAd75n+oXiNlIH/Io0+JuGlsUwJ8UsJ5j0rY5DWphpVARjTciMCrcS152/gKtq
r9lyhw5uzdyT7Avc4x6QGvgZK8BN92Xt2HpRF/8wDNFU+D3qJkYYxoulr/yb6cyM
jYSNbwBPgCxjPw9OMeA90M2YqRD6FE9fJrf5z6NkjNv4AYxoOxvXqHEc67kJ7es/
uf+fgBpuA7GvSn44DpASfnrmhCApQPCqddZEhYmOhjoiabMRXcQJWhg8ciMd77Os
wtreG5FsukobMiavfeXbYNbqtSAAJ3mGOIbhNJa18E4J9NoVgTb9S3Sus8TuC0g2
L7GbHA7kjnoxnFID0zkNgSPsCoo47aPZ8TQoid24GKERl3heMz3faf0gUwzsOMY1
3SDWKgrGM2yeo2EG/NIGkiccQECKwJbu6m9Uw5xSABJYw0a2Qi0N0YeyEjNRNmeD
VwHS5xo5y0m3c8d1CsUVs6TyaR7bxcaV1KfDMK5pfFSVzT30y7Ie1SlNWsosvaQx
Yc6Z3tCVx0S58zMFVpO5v4fXYhxjABUEw/pTtns/fI49zR8fXaSw17oH30gs886c
8ePbWNnO6GMXaR/HtYuVQiFb5D1HtYvEImHG612IEVUyUhD/UNyuwMLKFU8du2Nq
dRJQFJcsMeGAm8K3ODS04e5c7Q6KBvgIHxwa3lWXsEVjw2shaX747qrVKpdrWEMm
vIkwzSZdeeLfJgiv6Iq/7L/Imou90k68JgE1TDpTuk54d9Xn61ysfOapsGuuWCLt
2pPaXvQpLcyWMpo6qNNWGZIBpR5uDYHq6d2Ia4yDtLk39TWmyxEJdqW7UGMunJtw
AG3+AYf7DY9swHI6gRJs0wnfcakNKUYBkHbqPZNBnLR6cZtPsW14x+gB9JyHRwK3
v2/4mynwJboA8xfsWxqY4mUdQNCP2sZ6dzlKEA3V+3kEH/JkiXGmya+kPn3RQK3J
WUu0cAlX4YwsXfZOHm79AT5K2qLXkcQpEfzLfHbxNBYjUSuEt4Jwg0fG7nD7iSss
yrZOMGw078Zthhf5xraA94/cunPFn6on3XZXni7iE2KuCrpc8AAtMAUsUeGiKi9p
5z/kLIi073Vv3P4afoyFmL075R648UYmhPA3PA5OorgwrO16k6FHx5Lo6Ff7DtHO
UxTjRWRPFPZA/m4U2UP/j+ACtcj/clbcTr2XTZb4WUhzsEKrCuzNOLvab9rbPye8
QsVBcmRCJl1Gry7HJoUC+vLOtZE4E1I74ffw81XrwOsoG93K+El9FIzkorbXRaT+
7ko1uARxbfaLl/r6CwQtV61XTqfvrDdOykPUQkZK2viYMQ2WDbrRXXGSTtnXaHPz
YPCSsCmcOo7xedMWwVhtirIWlZSMB9bK2aWxY6M7h2r8xt+bKCdfgAiZvfeGwd/2
7zLWLAGs6win+P93It2EDQd7VyNxt8x8Rt7sJ2Jz8MgibYBLCWZg7jrL43AMlyE9
DZnk3FC+bPT7X6LaRtfcMVN06LaKuvRV0HolCeOYgVQDH/CzFSMIYAxxDqUN8j4X
tM77H4p7TwmsvOQRrPsB93ID6mYyQtjeZFwdOGfb1j0w8VLWa6qRtHYc+/XhWAPV
1wJqZwMfc8IVqe0V5zDRo6d7NGAszydUZ9rK4GNW5/xt8hgI6Qz6NpJuwUcHHhDi
5L7dTE9eF96lqapQo28U9fJADbs5dr5e9IULqp9orMU3opCtTzpu9mjCiGKtvjV4
5k/3nu7UxeUuytx9q3DCBUiGWaVMdNdD2ZmRPDRQu4b6Oh15CZkKb0ECwXEG4uSm
HpfuJX5owxw6WoX0iGIG/zPw38JHQ+Gi3Eb02PLOUJEQCiE2cOVEFRNZGcfjLema
d54cyj6bd78cMv3PS745a8o0DMrVvoTpi/FOzzvWqQrR1T48jczeUASFFviebrqA
F5utog3p4jBr+lFR4TOKwtPKHM6WHiCi8owEjixIQN8t/dr1NrH0wQPIAhgU7orW
FWv0GsA7FL9gKtU+nF8axTUt+Fq3ZmnZtBcKZrV3L7UQP4a44CoK5ske/9258Wb7
vFpadDCC1CIZm/+vKCGELdPk8VYDP9Spq5YqLw5g1VUQRyN+HHcsTzyAGrd4wrNS
3vP75JUrnwdvrwUObp8UVsHLLheQReo/cY9C8rR6KmKw2YuYsIDlgpvkzKbwPl5U
ajEyzfPjOXKXas4M2BEPqOj1Xxrrz4Vh3rHPwQskMRtUnTg0+E8z0PujMlY+KHTH
ATY82HORvIHhwe1Wt0DOY+WDsV4DHVnXHduLD4rV3h1MGvO6coDsLxHDz4YOQCwQ
MTecYIarFgl/FH+L4DAdxoCJvW+WznpAjgzpKGjIwNh8j2K9WoDQOR9GWiXWkHrD
PPpImbkzlKc//Ih9KtPeXaDCu9bp8fRjp+VJeGfGq/a0t5N2/hfvT41BKlhSfU0P
jIFd7mJXMw9gVSykOMEs7LpGQ05iuW/gE8bMBCZVMyYpLk2SSkU7XLs86jE4HEgO
nNpwanTazX+Rsv7C2/GGhVQecQVx/Vo4MyvVaPBefAgkAV1CcdxrOg9Hlt6fjpBP
6XubCKOqOw5rB56M227hqBjapt1+dBnu84xAZQBOkL3c8biodmPy0ENMWHugKe4r
TnUhHxQqjV7WCsmWboIyU0PCdmPkQepmJycF8CGyRZwdU6u1DSkq14WmSwLRhnUF
RKYxLz8r4JCkGnOilGnQrj7tdVwRo+Cwe1DjmbO3yQJlNZlWfHlQeGlfXbxUci9h
2fKd0DWRuh7SeyzH2AcYlqD/uqlKXIlM5rutBoCA0P5Hor/QAVjqzSzzBMzMH7la
ioP4/5Pfwtt3pcoc9Kcm74w1iTqtALx0L48JPi9fcA9SRu63WMFfzMEkePMTuhgk
32poJFmUKZpa3xAHDfIpEkHr1r9RvUbOmQWNwrzeFl+Pjn/m5nhwYNeX/mbJvKkb
tcmdIFTFbPp84PIC9H2aVH6UYrFyhDvI2vdDqK0yK3jhVuhKRci1d/Z1oP/XVWf4
ywq3eBiIMDSQ8WzVMkC0Ia9fU6b7gGtf6Tr0BQSdA1iNC3hmuYcaqTgxZbyEcuDW
wcYfWyQwYOiwMpPabp/le/PFgtaiEaXNGNk9aARL1m37FRts0j69G2BbpGVgRDKm
WhqLLbQrBD86rE95htN8/dvx8iw5NWQyoiaflhveTOfIEY2derbeAVYqv7lXlaH7
Ez23jij0IEER8/NT1UTcpQ0IKoS/0GJyCnbZk5MmXk5RVcXUjfQOmk0yasrrzK6s
TTF7WE/eGA6mEU7wwNoBEQzNsIjc2uthbNP3yp9kGZLqDC62ck3pLCOIj9rsj78E
dbZtoDFacqsIcuIEQVYa++ZcXcAqmyqGAzBgKuqgSph1Gwcp4iGDkMganeX7LNYh
Waf/eQNPHUI4jhFZN5oQ5vStKQo3X1TcdgnHZZFDRkRgP6LNLpIBqBqYMdFA+VR2
BE1+aGZp31kPCUWFqp2dGsVP/Ai9hUCpgBW9aVXk9A4pdPqf9mXZCsnVFMUVz1DR
lsaFvaM6Xz5qKisb2Kc1qdYcu5t/QCqn/Nokw2PulfWKcyrRFrXtHP3Xdm90wKen
1Pi21fPiuXOBUBNHSOm0SdtX7GOOaq7VtBlKhgYWuDSnc5SfIPrSnzOtBJg0QeTL
wRugMJ8RhYIPh3wIoxTzUQvRht451XaQmKSeaYO7ir/AmDhdQqZ5760OZ80gunJa
SyVLJHoXUSBq4m5hnNx6Hziukyg+WV/SaLRIEsAbXMN9sjoSLRbqgSVJXt/mv+th
ghmDhkHR6spkETvL6gdrMiKgycq1WAHvObN98basCtBXOsyi8KJAy0UGMNpjiHEK
O81E7DisbvRs1CW1XERv4wJznryiSc7RUK9kIPNzPSYUoGnGMbVS6El7PphzsFh+
g7FVU/CodwKyv0cEYdYv6aykXbG/SmJ+x6juo0F/nweX3LyyPhVxKkHXilZB59op
UGee5/q30keXAWOagSHg9YSzZ4ALA3Al7iopT/IAXRZN6HUm3P6NiwhB96XzlJA9
Wq+B2lQJ+TjtgCuCFBwn+DvoZU/Eh8G/EVumjG4lIQUH4LUqlfl9VZQqdMzv0/cM
J6WvsiTm3AtLTQSl5WG5Q51arGbMIC4y22FYSsm9cD7dayvW2Na+9uvlrnwvzSRE
zqKtZ73VYuj1uMXoic5I8tMYqllKrA3q4E4lnv71NZOlR2cGjSNFnTrHlwpRKSnP
l1Gx6wKmlNU43Tjx+n1kcD8gUbOpGcwP+xQ0C8MGLoAO5+KbJWcHe6EEdM0ja+Yz
aeNsaCsfDTy12GS9LyYBp22vTOudTfnZbVpxvwSxgOdux/jmaCZoxTBF5C6dZ0Gk
8ax+rOMFMUat4fu5lVOV+ADBMzqvOLZFrBBMEfO00LTucVIv9M0xRrdy9mkpfEvR
5rQBiMUVa1T1mgPcvWs9tci7FIfwYJmVAFlax8tYYc/6zbLgVs8r+nzSZB+cS1r+
eQHPIstMrrj/qZA0w5wNH2YpUEXWET4V4l0dO0VQectGwVp1xled4gZLN5zJStvW
l875sJmKKDQ6qNwaqwk0qqKt8Z9tQWpHF6JwSd9WAG+2qqfYuJW02dcaIcxe3FFO
dWZwRS/peeaE+/3AeHmlzfwLuCjc1qkgWDCEbq3SCr21sdFmd0mG/kGC1TXKWWSX
3NmXKwRKrGw+8mPDKxzyDQEXmAf2hDwUDd/a4TeU91NH3k3agBVNsgnhyRsC3NVW
8L99WPpykBJh6mnEYuolDtCMLo8T89vN64RAgs/CdL43uneQWExUYdsIt0nPnfMP
R4lA4stiw9nHqYN2oExJATvJ4mRmHxfQO1egPkYV33BRWA2TWScWbEnHmffgwcJ4
ZvQmr6+sMGzA2RqNTU2Vwmksm5htxvHyyz+p6rMhOR3enXza9MlECQ0jNTDxPx0z
byiIHWvZNEZNDmuqGo5c2QDiP2jlGE81JqgfAkHiPB/9VD/zFKYmdBMfsq4rzOGX
53Io9ix8mRWijg9l/shYD3ziEcIC6jZGSDPAp1dxTMLmE3mqusxXgFSJ6jm3tUCj
MGd8TQedHZsLlC4q8CpiOZNgwwA5G5eqSEVpfafPpGezQ3FMjdcBvZZemB3SJ8HL
kKeehXvQ9h8AFV75k7t0pRASzgZAY9yTJchgOY9FmEOixliBL3m9vUiCQ58BVBVB
sE9yso7x8qDE6RkXh86wF/k43L0WklCRucUqAnSDUJDTeRdvenBQvWq7dtTTOMNI
eXlRYTv10NumylsSY0b/CzflbLeOduy2SymSG7uYxso/yXY5e8dqeaGeNHWQpbyp
rsd28g50LUSO5+80+IZDHX9dGfzhQ5CDjPeR5/4SVYblOfuYT0f+XXiH5DRiNJCG
Nf77bqXV8UM/j1a0Mgt9rgsI/QBK2OHZ20zgS7d+wuXU3c9rEibo1A4sGEiK4WnV
26XighjeQMHqJ5PqzqFFJIkG+rtoSkAWf//ZLe5GdmijDyFR5Ky0UMYl639KxIbt
ozke/OiTnYkTmIGSQOPCPG3TdgfLaHYwSVPZF6sH0tPJ1KbV/HY/4nzv5MXPXItB
ou8Dmj6SiK0KdatZqLrkVceDVT8iPtulkqbF8K2n0xQJIddweTtlnGwCNCiwNysL
pVjZKSkqu/cIa18J0O7xc0tD7aPL06Y+e0LNJGniVL9wyhc9M8skG7FInA2RSG4q
UZlEDysfjNmA4sKeUwOMzh/lxySddqRqfGb7y1R/sgbFzZNDqKEH4cnp6BcQdMCF
i6M10Ose7u3yao7/qqBtvHq2iVN7EzhrIfL2WqaAaeMAWbr9LuHskHZZqC4GR6FB
0Wv9oqKt6bA1h9ashPfhdZIetTtPI8mKzX+7cPwyO1cNfB1B428oV8g6CVojyy2/
vkMWVFKh9x0ppiUJ1EGobQahugPUSm1eBJ2iuya+TNg42c9ztvenrL6uN7pnPnJR
ZmTUUt2qCpsMcl7OTLCrMkbE4e1eGvEUb9A8xNdKXSnIcc8ioOtHFVNlwt9COBr6
ysJz/Uuz6dqiILZJ8p9xLYA9aR2LlzFRlsujFWrZWvsBtkg1jdnUExjw0MPCPsU9
oO9khSBBYyuySWdNSsD6DrhuHcd79V3MlpqXgjFOpCQfpEFbvzhQJYf1HyNuv/CL
o8s32AGeiyK3E3JfmJyFMIUsuMG3sFbgcNJ9qIeHWMSHyqWc+H8Y6AwRMd5bBNsq
9cOSEa9JKuRyNM9lvSfAavxY6rRXc0o7fy8QjsF9ZhT4bz379iMYN+wto6lCqbkD
RIHU25EuFcbf7x7jkHTH/45oaQkesO9P0sQmrGgyRqp3spZGnmiRY+4Ngcq9Iu1k
CahflXKOG+nmm/xz1N0BLc+o/o13HE6eqKMdKRYRwUagmQvCLtZxZn8axNdlMbJk
eZlsl8UQsUXl/4VR4CCBO2kCY9DUo/lygHKJeU3WG8e74CTVKW5B3NsY9AmG5Wkr
8AqP5SVpIaUiFcniKOIrCFkHA8WVntJf35NWlZQnoXV3WOuZ7tl/90U9iI1AsWSu
oly2cT6mJPDp0ef/oZApuv1Uxmm8EgcR50GIKiM2T8pYBVqwRKRBmL+ppXhZbAZf
ztpFoESQOHIAwgOZy3VGySWvRJMbPlIHJV2DAkfXFuUesW5vSKZxL3o7pmuW6sBN
2lU9dP2HAa5roVM6UE9ur/7CezxcAU20A4i/DTRe8OjBAEA/eLryWcU6bI/5Qvxi
8/fGlxbmqHS3MnG1j3raBioFJ+nVGrhQNqGHmwautEM=
`pragma protect end_protected
