module crazy(input logic a, input logic b, output logic c);

assign c = a;
assign c = b;

endmodule
