-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AWOkfbKOa3ni9Okzoo/Wp1saK9C1MFj5vaSJ5yOQHwFhvi1Sy/HtKufJ3JwBRKQJ0jJ3NVmgU1ww
9Td7Pe+G7loIq+UjV4wR2aqLnzOutHOwVbj4rtCOMyhAqMWqkbdCe+XXn6NiLbi3CvUMf2BU/uE1
u48eTiZhBQzHaakcvrTm4ah7FvPruMUmZjASK86ExImNWtrRFCu8c6N3br8Yg0nz5U+4pkR5q9mJ
N7ENjHLAz47SPPHu4upyslCv9lGRLDGcju+RVMgTpLsVaQqCk/O4WvpavXXSefuVrjjFjeKMUcBx
A8Fmjhp6SXOezzR0MgewI+9Vxiq9rjsom93r4Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6672)
`protect data_block
eem8yyH/SHweGRjK1RvceXvwB5rGooJPYdgLZqFs8Y5kaaMjdIBntanIs9jVEY4Jr5Ya8L9JTCoM
/XIdimjQn7yM8dKrZzzDazPnmAk1tl7nzIUpX4cKTFLFeNC2Y8ppK0wZKWN64qCSvnO2K66LS/aN
IlP5myXBUMVZ5+bnGMaSd4kAiAbo/SgLmJeCzKT2CrwbKLz7CctVREaSWI/8Vb+kzH1kORjPiLGm
GXPJZqY+/ZeMxRbysU4J/1SMzpA3aGnA6BNcSRXWVZNrpZB7HM2CreCjpzg6Rz79SsIB4KfJ8xgy
hBxeEJ9azVpnCiEAmWstq6j5z5gBiBZKLYnuOhqJ4Tz9nb/ReVy+RQYKt+zx7bfCpPF1wxDSgkte
ATElFBgZ4/NjOpt/dzH90IeNGQKlXLXyzrCegGSl5pt7rtZRlFzgLI+8owYrooqQdpdyZ76D9KTV
0nk8FTha8hsvv3fQLIvu9yi9ZdD0LnBFI5AVOjMf4d7BjwtaUptyVVV6u4nhayEUTwvfpYBgAaQ0
pe/YT7E8rArx6fQx3VI9Epb+ZKCFhWunEnwvmC+MW3VESU7LXUVwKhTu1HBneKvvvMSH9wCLSf6d
hWfkwd33cG4PpFutbdgMygWqMhJMyDz01RPz/4+HSuM+TPacgW3/tuC4ctfpQrP93k70rAZ70AaR
xRMBhnsbpOI0rCwoldMtA1JXujoDA1cFffcZZBbnwqlW1iewIE49ngLPd1zCmZlsBikma3sGD3Oe
Ov1bFnYErnNJnpMQJusGgXhR+P6/fFfhln9EZIzVJpoJ69hDhFJi6n6qco51cgCwwoPYsAVv0YMG
BuePlIKJhjrW8cRNocLDtmlGEhxwf8PFFeWjN91R28M3Wg6zLR/GAQWJoLAJEhDWMiKH2dGGr6mE
nVaT0h5n4xTIhkvZz5gNN42F5dn+xF5241n3J33lzrQG3bwCXcdSyJLO/7ZXwsQCe5ReYUdrywwn
R7MyIqi+RiaKJPY4dK44IJg/NZ94VKKiNCzSndFIYgfFKWgx2vDzbafKf8zuaSuN6XBQnRw4226E
aCaf1uatvkT9ZAD6xHxhITXYWVCJ0TBISZ/HRXvUvzzrd+dHqzeFUNG5TSvFxv4L+ULCSVJPwMcY
NvqWsunSX5TH7vyHep1kCCweDf4/VLv1XS8H5yKUpcJZ9EPzX/l+0NFuBSn9HmLZCVTawPwVJVYw
goefy2P0R0pGi9sY584gEmBNBSJNRy80InYoTI/4oGRx9HaZ9ipDCvxq4BkIu9j6zsvQY8SbCU5H
ljxA4SDCTYl6yBYdGYSd6I0rJ33Zh7EEE1d8jg4w2Ur0kjrKsUv8Tj4zwE8CfoxJVDDujMXNM//0
3mK9LkHitWqR8GWU5JWYInoL1UpjhVjFOeoJirnrFQOaKnSzC8LbJP9w88Tp9+Gkh9xo17PkXqcG
UBRn7pj+4xdAZBFjRrEtEzWwJPF89ddqdvbmZIwosoQb6mFaFPZKKjtERbbSSHiFBpvvWCJwqSwS
8d356/A/sGrzxZwRxN7KDU+hU2IjGx++O5jGxN2ZYiPH0tqGJnFgFH9txXF8UoZZYMEYuy6aIu3M
QmML602Sy8gYTMX4yzKwVN0IEqJouQWgLSV46mMB00ky+tJFV66vDRO9lJylFTW6EkZYn8XKXv1z
H+dg7jKgLQykiwD8IGa0jSPW0JdBBrVMq3cgvqSF2MB8iyN6Uaq1Nmgl7zY7cQslhQRKeY3cEDL9
Zjm6A+mFdasspdfROVID/mQAVS1efMZZkScX4Kfe/gBoJ0k9EYt1VgOXwPnrqNbQ5A4DIaGw9FDy
O4nHAt0zyh2SKXmkC0vchXYs1UkMeJhHr7sop4ny6TMSDY7GNTNgONmd6qnAVHAOzoaU82CtW7PC
DWlL45bO/cRO7rXjrdbxyjz0Chbfr5PnTR5eVBCo7+Ylqa6lk41RSBEObL2c2bop++Pe829KEIWs
iQLHExco/7SgjamQqKIeqX1DuljrTdzl/SbzV7STMtSAKxfL65MbMUhV8OpEWSGNvRbInkUA6A5N
gdGJiPgDtBYFVLAyWQXgzPEMQ5nVgMLZNcY4YMiM8RM9eretFWfMaRKNqvAxzDqv+sP7tQv/HQFj
ER12usGrFWZkS+W9rMOJm+7Lg6zD0NIf/VnM67/6R7D4y02mB/l6W7egEzUM8Ua4neLFCsAXMtZP
pgJGOAl7xCkXGHKtMvYcrp4Of7dkZIqJuEawPkXkwcd4u/wkMhykYUv941a5KZTUq/zbOirz05Kn
RvrrrIu5Zx6RwTt/WgLKjdgIC/QSoJYy9yukLgw09V/fk1M4F/XrNcqcfGbk/rTQbDLJj5JBpO4F
8ZJfnn4jpOjcQe4clvndFYqltFUIjR8SkxLaE7jV8GacmYrw+Wh7Ta+/ZRlGgnhA+zGQMeGMPWhM
V5sbBjlNu70ngPgYiB+gM8X5vbtyXaqibsngMk8zxntIaehGPzmd4iBg1WM3v8/PpyLdWIitvB/o
7oVHGrIp5JY1PWQM72mN7aZZl1b4XjQ6n7DJ3gGnY2teH1EWk7m6dFa+F6qxOg2kJe6K+MARqCsl
wy+Fp6YcEvmT4ds6yUv9HyQIMA1z+xjKWPddo1109ee4fteDWs4p3JsemT+PNolVAEI9uNpPTyGb
y29utIGab9luvQRISH2+edRWhPw6baNTiG8roUX6oJgOlYvqItgKDMdM6sis0jJg9wlKCLogCU47
6ezZ2UbevOpsgc1CflqnoxiNRY0rRKp4LPL+hA46EdXnHbuIiM97RGE99/+zEjlWKvdFMPnxO4jr
zovyBU02+ImJp1LO0+oXPNE9IaeT0i1o2bsz8b7TUwQS+yAOGTcQfYpiHgmf2T3rrxdTnfH5MH6f
QSZKbc6iKmoRMC1b12pe40eXWuYcRpqtzdwsc2xaerpnFPPd08EtpgFJhXeTfiyqIYznhjRv7LiK
OotX2PelMMqesioYNLzSMqh3bt/bwNZsnsGgAjMZVX3SOlRjX1C4t/ZSG1RILV8B2GFprxDzNck9
EznB+op0WcvTLilPSDhjuuabYZFMcncMK+uk+h9YrEqaGef1kx1Vy7Wl2HV/kFU/oh7vilEOjU2e
ubB9J/3IXq6Ptlw6Gy+D3CU8qfEJI2bKoDtSbvYYSGLMSy9Q2A+2P3SRPoRVSlkooxsA9x4hi2tC
YpreyJy2gG37Ym5tnmWJqm+CXwSictuqwyVru/mwlNDT+KPgWmbRuVnXXVCPA4Dl39wm2LtJSbs1
ZUTdomXcsT+HtRwErXdVt1VxTQ0zx0RxS8TXy6O3+gWVHDDfBV3xHOT9A1BBf8znD0Z//9e1szQM
GuvQhghvKNCZ3VcbCjrzvzatyBWyu0x7rHnWtyXq3FQUDPyoMBrbdbXbh4aF6ejWkhBvvc+S9Omf
VerZflNPlzZC3BkmaT3DjeIBYoK72Nt5xBoegXz+yBKsoLu4fXeWa8/9Ue3OYFr6he85WnzAwzYS
cyZhnvFY4r62ceJ5HJGyQBFTg0gKX6sM8GbC64WXADdWHgc8f2w7PX/qSLdLq41bOnZLlWyU/LZL
I4AOVX+jsYDfO8yMECiWhEWc2j4wsQ38Avwhk9CsXQ7DPYyy6jCsXvt+BRTMmG2zKpWFZPwTckQQ
Qp3RWJvU7YRo9+Z4FMY6ykOgDy+63QJ3Xk2sLyG9bRKcBrpZIjMqO3PvRq06MGOWrn2nVpLhm7Gx
DS7dE1+EXNLP76DldWE0jKBneT+AiZA08zg05cBlmEqMgdfxG1CI42P3qPgqOIPlWgjl4yhFKpoi
uG3Z/HIsO+5ucbJcyzBkIh05ijllSQ14AWoxqCy3ls+JZhglWKYJVRDkfwtqqUWPfPdfL69r419b
vx+gOcxzrmsWC6LQZ+vqDGPgNuzlCb6l6VDqfORJwQp3uh+r44CXIXsRejSwPA4nK7xAh/XWa2W0
GDWksWnQWyxTRAwQ4Kb1EbeyI48t1HzVEFAANN7WejIOk7230Y14DchheQSNGPjVpowF//rYOAp4
gx469BZ1LuApxvCK4dlnpEjUqeSQ3PsdPc2pe7hLWtXJenhhKDKvPI+PUFefmzZ/SsK1mCmIftYY
2GC5E7i7YL8bUFstLtT1W7B2Y2qNy25Y7nBLSgXwDW/2Y1VQEWz/t2u9M1s2SGG66N0cX9pRFY2U
SZzvn5D9T5IPl6lbqQfVlyYDIdLk46+RbJ+Ahs0w7V0WKefNnnCbUzXV/0xuh6TQd63rvssNjgmP
wbGG2cHSxCdl1Y+jKLOKL/s5mXwTRSF0TQSANTnnMY63asTxBNckH7mNs8gBOccnkobS2zrKw1bd
jQweZAnG/wdTMZNMyJl3BOdFd+UH1n70P55SO20SvOrlVxVexdSpPqHIwEfQqhS0J3RRNXkNddpA
4k5+bEFcuPHtO1F/OfqqTs1NPPEyOQG3sgsSLI75D6mQ1OLvyDB1AajbLfzbRfmjF944RCt151jm
3kUdPE4Xsuw/OtoHJXm9nx+pnrbl+NzKnso0gNjpUIeI6gielCENkq4h3YcdLM04KwYI4GQuLbzc
4q20KY/EjEY1ZmIzkbzV6u/EUSG3F6hRs9DIlrBli/MKhXB5ABdhXsITg3a0bTAyHr6HSaxXDmxg
xl6ZrEaMWbTIEpa/xiAqkfFFCiRYHjZbdd03HpzrJtRnmta/mX4vQzaFzgYiJHhV2AR5RrVGA74Q
inayYBImHuXWP0Xhah9e0pJV4WRgbWDjrL1HMvRPdW3TbfexHghLQeGGNqSknyT9ba3q2RkSnHQL
ffhn6c8qTzwZ2PHldsm+ygbSQjriMdThSqWaqqiurfWlXjbYHbxs4uTt7qg75/SpU8Ijze0YT8sU
zzjZzQc4qKmLEiqfazSJVmYptMeker0tntSrExuUTX+fXYMNDtiBz/VjbOfYYecXbiw+sTvEeEmh
0qLnPtInkWk6Z2JAPBnB14PKfB6eoHzbLnM/RZDz/YdlQpQPfjUZKZKVq1MyyKGnC6i0eMbyHsd9
O/Xu9ofTorWRQ0N8KEng82Q8UFlvjSXScha+MU0nuKyGXg0fsshTpYYOdbAQswdmwtRF049vqCwr
ZYEbMlrkwEh5kWDplQ8GMxf+eyt3Ir+xLvr+nMjXfRD2iFE/lN6t0lQkcQOzS9itYRpvoKf66eEq
6NK/o0fGkfeHMVtacZ5A7eIRkichgLwaM9RId3YlmISRQdTLqnEpu8GCMxRPAoUtuRUUl0NrIyTf
YbO/1ycx3sYMaJF3EyNTB9Jzwue61D+HCEtDwqSHfjcBW7pxDtOw5DaARB4wtWsGAyMQSOCwQ9iv
+9oS16ayckcMXh3zSC9KRbrPaS57Gb8V/AOxttLl5X9QJW5nbPMDxHD0IJO3hy3nJ1oiaVM0hwDh
cR6CO6p5qzkTyMMfjFWc95/8t7ejWmEStOkkKYmVmYPb0VWAWlISRHQdq37d7674QGK7ihLwU0ie
qqttVr1gMnmr7FtJ9ygFJGXT2/G0ra8xhwAwLNREXLiVPVSCLcUkwdpq/TdMtLgHQhh9xEg3dHlz
C4dp5w+Cwh5N3LjAUKL7RhQMmrEFWW63qcnfPYABHjnZ3kIEgWwSyGncgyB33T9VlnRLMgZkn605
H2O6/UMNd2whS3TRgS0OMte4Bw71vDCTqy1a+51VGgEqOvplwIbMxGwW9T09QEn03KSFv6aKGC27
dZOdfCJjuqwh7OCe++frdW3Cks8IkCiEv9Zn0Se3QE138RSzjzgrDG3HI+FNafrFpXPwbIJbr2Mi
E7uoSwljPFBlJl0ZWkZsvrq4ibey9DdkXGnOMouiGn7uF75/nLAluQIP0RNes0nrpdiEpLyBuRQv
Ff9e5M5OzD6ACmVcY3BY9foB50qM0k/E7gVr1DOvyqeb/jC20n4mm8tlweNsnLLU0fuxXkZyXSnd
be0q0OMPInATTX+EVjz0sRsKAaSbnw/Ag95ky3Xwy2yTzgzG/lly/BEZLGe+kOPjYtPVJib/ygSG
3qwbG6VxQWZUWW3w9arhCLVYvL1ApkfCAV2S4TvgC5wkDm7+0VsydKn/ZWhejUFDWUUfM7bgRnAG
a5NuMbRhaUeR8/tCbIImp7g3c1WMl4wmnAUazhpREua3HTld/t2lmxBpCB7fbmtUQbEuhPYVl1I+
GZx9oIersWanT6j7TyOZjeQZa2Lm6+nNmBjSCslXHJsm5IEeXo6v9EDYDn/9uqpEoJojxbY+Hfey
GpgVzxa4sNaH5mdvlFQxbV41RMyg6HmCvIiUzohbxbC0wMTS2f1aVrXFIsu9O4Hqk7TIFgE3hggC
R0voVC7ktfIP+u/hkn+CVWGVbiEceSeCcojHj2urWrBRe3pz//wD96aQOzwmQz1SZr/bWktXbQnk
D1ndso7uOWoRsc8i3d8epnWtf/L/XKDNquOutx+LfxXKtaWh1lDn9rtHWI4PzdS4HZfV+4U7uS7t
3RfkcaD4DG72dB2Xzg8R4zekiuOEpbeEcoPQZzjTHKw0EZnLlxtLyZ59aJr38vUWJefUTqkGLw6R
Cag15nkxnicRGtDmZXMZz4cWITBE0tnQMkC0RmB1bXpblvr3hsMSVw0WqMP5rtXr9F3W96JPlmqy
1DBuii5rXU6v9J6CYl9D03G4eK7SydKAV0T8X/HwmHG9bcP9hASLN7sQ0GobRiH014sctbZ+Udhj
nWvvSoNk+9FdIGUoW3kTNXJZfWpw/5BmCbd3cCC8PjfMPWdEO9jfVhOpBBGBdWIuYVP3AyTOMbLx
Qg5CxfPPxJ5yJYUX41v9ela2d0tpuJoTkeqNAENRu0wE2GIKYNs3Ks8ofMfZwfhS/xd+a6OT6KqC
B9ClyNHTUt5rWglUyY6eEmIMKGdiR0dn2LfU8xI9IAlNPzU2pikhEcnenhLizJ1QSBD4qNxJGopa
51iAu5kUAQ9bgMsNn7Ok3JzgUkenoKa06F6pFE2P2TOFEeXXx3xA2U4Zbmf/YGyuaBr9rr1IyioX
GRcG5VWZTTV11q48fz/RJOUJFjIJDE9Fkg/2MNduJh3Vdk0LTFpwDAvz9nTV3u6vEcHROyoaAMCf
qfyA3cJJLyVLYgQbMnNPC5sNSSqq1VUY0TIZKEH/wtpwNwDK1Hu5BJ6CRJfUc3O5ozgkS0kt4Zsj
vfhBdnenONJPNe7dSvX4YRufqs0HejItlO1ZwgB6dE5VDXH7IQn3egcoGGw3nl+61KJ18W0ekVkw
j0IHCgOPFWlCUEtGAvXaQts7MEHbVLlH+irQ1n4MCBmtlEY876cTTeeBEpGF04bJxVmVAu9Jh9mc
FyKj9+nO7CIkhzI/9kEFcmMgMgCnrVffbgS4XY80O+v7eFR+gd39Cjd2mjbSz/kCNw/QDBga03T/
tWSReB+/w7gBpIii7A9hv814eCzR/ouxctsWvK6FRKAZj+GoTHEUOQekw6N9ni/4MZY2vuU1jIuU
FF8drdiXmWJGaKHNXNhaHtMboBS50za1fEIN8pY1s4YXiWOokoPSpndpDuF3MxjYVjfC4lfOAFF+
LaQqGXx5OS0Q9sgNxU+yP/9XWrFlFzGmJ2A5W6iA6mh6PZYuDkLnLfFc3xreXDDZ6l2mZi3W2O0F
nctd1VteWM+J0JiDcYBY24BGBBRbGt9gvvIPdEU2qtT5zU2sFpZF88YIx64nvz7WDztbkeZXxPtd
vb/RcWfKexQpbeCn8rAcUEIZJE7lNx51anNvPn4JfvrPHEnUcbJ70wSmv/Zl9/O26s+W6qDBH7OH
lze1DIby/hL3H+fJ2jxneL/Vm4LPZ36f2G3ILUqKugGfs1yGlRePfVOGpusMuX0NQdyu54d0+2d8
2tWp/5S4FXqcvay2D6PIr9C3AYzetyXMpJ4XrJjiXe+Qek+9gpVfZ9zXDhTbn2e+WjNA928li93a
pkJO074D4vjEdmcDeQVW+m5UD4Dbj7fOcyEhn/+t31rw1UExCy/dKFoNyS13xZWrY59/8VIdWYN3
jKnvkHlLL5hYnLIBLgU4QRNnxz/E/PuC/ZY5HU1aXpTHuXkXw44vqJIjOFLycX5dLJOc7E2EXKgU
jYNkZWK5Znb3s76mQtjzk00HD6YMcOYY7k89dpGs6xkjvUrwqQTjaVkPQoS4QbJWQE6abSUVSPxV
xqCEhdvjYXUIXOBOa5jyryhkiREDN6fU0j7+NjHTdzVipzDWMJ+NYZ1kBq4AlzXjnw8NLPELGCgw
mzRMYHjTzaqXZD7xD/479RXSDxVVpIKvJsxjxlDJZq7HP4MpWxjdTFhVi5ZiVkehLwa8ykfJUnqH
wZ0WL543e3qbbj3cbXn08sHGxri/feidrNPLwb1mZuXDyHjCCDhgZ1ZA++qMMBFUKK4QNAY/hKcp
Rk1kcwI9wym4waR2H9+7oUEk2qeNda+a6MSPVqh+lwLVaeyrCU+z0m9yxn9xa6n+eos2oiSqNS5y
NQpR979bv5TrQa0bDt5KKEwEAHHbBoKEYFH10OmuLZRxFll/I/naKCaxhDMadgpfGYjb5aKxHji9
s3kbMvMiaXmM6Ici14UeEbc5QhaD7y9Vf9UKW5B4fcBBPgusuzOgi03rcxM4NrNGNuwiPAZIhP6Q
6RGf0Tg10WaxEmuqhLLuDNEz42+WndbC9Y7K2Gk7EjukJDxuCRXL4egt+dIhwFTwylqXDDPYK+YW
SvL3A91OhX1JwlI4kVR1NgownxvCDlOcLz8/jTJtLdXTc36n8kudDVeZAG5k5wVna5eNmtIdXJV4
tAbvUbqG4VMM3nLlYPU/5gWVDis8kp5og4peEB9rn6xT2UUOqa5lEvSNTv/4pLmzXaGEUuhVjt6C
poNxo90+Dt7zeznOsCsxVZRofBZeyEWtZcmginurI8lfuNkZDx4RirInXYTP2P1WPrkuILkGX5Ox
007J
`protect end_protected
