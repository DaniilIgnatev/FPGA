-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
x2ifidsp9QuqBdhiTeCBiWHajO9nwbo8PvqpZuwSld8ALCcP7RUp4tHqSRFxixr+yHMdJtpacOn8
nxfKklT/8cJDGX4BUk34Yx6LfeB+2aKNiTcHG2/Xi3owXEjyKTw5OshCvcAGvhCupYwsA8lwXDWG
dPHbeOGMpKm3pkL82HIyKu+8JNm8upeH5YuuzZz+A1tHPMdsGIuQjSdfbMZlfj5c6lhC6puT3Ygy
JcQHGqV51j68Yh1shthdedIQq3BCx1qu0LmX2XXZ9I7HYPT4jm4fqQ22VWLSTJjzr+KyglbwukpJ
X3XPQpS1yunCEQwZFfySMIvUdU44QrdhdxMC6A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5328)
`protect data_block
8rE30ryf3hciB9eA3t+Me566y0cMISAIRHT5AqS0PXviQftO+Xrv9rO6h1615pRfrRdl8llUvmEa
lQ9qooaED8Z9kkyqX3YxMiHL0OBIgkU++NE7aIgUWmPNwfXHWeUR5ZCDkj8AFQK8NFUN//UNT8Vs
34SQP2H75VqDIu2bVQ2iZ7VQikBM9LoXDCO1yvj2Dva6l9W2mZOoJXieTY8EiON6UswK10O89BRv
XoNPlBNNmVXTQ7zfwjHSP9iH4UaQ1WAWyuCzW5kJuGk5hE08uic5GF3VfA/GMglB17ZDA/Ls+OmL
6SRf4pKfEtqEM9LJ6X0v8GPCr8oMLmA5JgHJm2tuZOJVTw3wPORf3AMdABKHmNwGxYxP0grEM21P
Hm9AN7OCFuwfxJ5uFmGfudlLaDGQ98K/fJWTi6uO0V5aTN1VNxbMzgVreQrfgijtm64f7SM/zn04
nXQN2nU3qzmqFber0yPiRAFWheeGPM5+zbTriiJkFG2iRscUrrwnPJ6kM6o9WRavPJv4tiLJWI4a
/9qKVGlU5A3KiZQ5JcsL8QcZgCRI3UHvBzuKstTPw1QE8oPX97Ryofp6gTOxtyxSVButNqhkMLNc
AX0YRWRoWRhCrfRNe686GY1CF0qHsx4ae6COdgvXcXArMiNx9th6KqmKINi9nrAcYH9HL8wbZnQA
Z9+01uCRwgbVuXH0EuES1ktdf+myMXHe2v5iK2FaRkHnhCdlMEusuSBccrCDzgEWP/qp6hsTTb4n
/gJmIhfsl3d6yQN9wQY2UxZ49oghgb9w9dXiN5+DtXcPf6Tb1HipoVjz/6qzYIlp3ok4wg2fCb7K
1KGlfQF44tGw8kVWVsOpRS0OQ6BDeZKgGmizWA77HCyCOK5vSzm/5WZn+r7Dkq8/nT0SHQ7mU9M+
UPIdkkt5d/ea5J9/ZUPvIs/aETtpWawJ8IK1a4qV0KJx2vJgZh+MuAjEUKAfvnWr/yhizRWXiGNV
+2l5HvdsZImdBIo7bVTclZOHxQ9ex5KpS8wa5t5W0N3xVRpcPCoBFtj58r82Nm77RAm54SnbTBLi
RJWfVpCyaioKr/0mkfh3ZTKpDs+Tsx7noU8r9cMj/w+cVhgbxfCRSnHnlxhpkNdeYwx++DuRSShU
rYAgESUP0/k0LRoeckljtd6jX73R+xiHfjjtl8hFYgQbbA14eO3U2phfGo1fFsn8AsrI9j9D+SZ8
WGczvsHVet3poq+crTaCsLTUMB4iWx6TFzGb5n1i/nohXqd73drqbhsEMPnVv/5s1NBnq50bouPw
PFS6owm+RZ/3QYR5dY8ynA7mJ5Z0SRtYkoXC5gWSsvCRgw97g1tQJBe0xHQTPuczq0QLZf/1IciZ
J1/0pUib8ov2GSxenOG3kLVjrhjLvgHlJv7Hb0sRcRy1d3n/gxrvn5avUmZUB1I541fOrGZ9DFqT
qIt4wp0+7qQAh6GNy2qoCe5QETjhzyR9oJg6bGveuqBQWGMVGAzKvI+drMfROZWRDAIAd19+suhb
VBYqbhhXO3bbwr5z5ooLfAJ0om9SDTvtW/vSbzr28C2l9sZMlZDGGbryWnVbXXT7KfziW/UrTNf+
VsxeavkWjTyvA1PfwHDBGQVwLTvnLdVJ3NWogBYA3C9TFj/FsIDHXloZRubld8J+8tyFZviOzZTC
VE1TV+ZECvMPDXALqrFIvy+4fcBQuuviPX0it92TbdMVIzTpzHEmOkUCh+uwODGHK05+SLIP7b3G
Hfm8WpMmP/QEFeEVaLpJECYBuE4ndYRfsSa2fBC4LAXT/Ia3+zg7xHdL6j+Z0ccBhL3Pgbig4jv7
YfPAIyMxuB5wX43JsZ9KvIQAbeZq1fM+nDHriUoeEyWk03HT2JY8ptimfIX9HX33+1QphoztJg9u
x5m1U3sGEZtTkKTsZ/FaChOQuzelMvG/ssXRjY3QtvGyViXuPhBbG07eVhcS2/ygaGAD7tH9/m83
vYSxcT/X+Q0G7ABqMubBk9p6/zoUCIBQZ1jYIKCdQ01KPvm3i+l7+9TilhZ3acuLs21H80EQ/ci/
JykCZU1a/pYkfJpFw0vyCXPv+bBUMiaogqxo3/2LkQ8P4FxGRUpWOOC1tvCl3EADJHDPsdpntcfJ
MqnLN8rmcUMIoAZu22qYOhzn2y4IpznkfGYlAeqyIL7uuokhpWDPZHMpNFMyxlM0L0akwsPyyHeo
fGkGGJUrh8gYlr3xS5tXsnxVgFIpTbmJ0Q7CCeh+p+nrgsbTma1kYrzHhdHNUKgsihMEX2JaGxVx
Udbyl6/bGPxxXrtiuBifCXhK9jixqvUj7+ICeDThq94WCJSt9ZFcWArLOZYZ498MBWLOxETWBgbj
ixZqJhqJAUQcFRXgIoqVmsnXIZaxqu9DEo43XEO3g/N4OLS8YXccQ7SV865c+7I2Nys6dVgMf6Bq
fyFCAIHXuoFcmVJvxszZmsk3GKKidPXgRi6fKiTZqGUUr3sbIXpdK5XjYLhiTHkr42loTzxlGv6K
T+g+5kMNppE+x1WUb0DjN/zD6gRfOcuWXXrr0BkiIokljtekPDWD66SxexMoQuYuYJ8HAI1Vm15P
zU1p6aNvjYlX1GDMa/9nhNt6TUx6f1K1UNU0AwEi8rvlBkOdtQMgJQ5x7FufjbRGjAxkUmYNwfh2
fLF8M3pkOX4zAcerS2fNu+1zCNUDPl4EzWCkPQ46WYpXQeZV2j+R7T/Fdwjy72hOABrLsnQGVX4e
AsPXECvjJeqdSxEdU7engT40+TEwcVYTFgF71X0qYG/Y0r6ZO+lxkZPAye04oyZeBAOMtdyTtaVR
D8Z2x+QWdS7RkwEdQphh1SLIDqNlRxY63ITW/WzDk6xqsMvXGyjh+O53+TH6POKWYKJWkLzjtge6
rajscU3k1zE9Da7+K12nAk6SlWBG9O5ySGtCIWtOpjckUNajqct1J5xD9lYVVMx0x7ligHvE5SO3
Z/PkA7PopMG/nnU2lLXBcakziNDDWJR05eVYYkhp5mg2woQ1BFgeOLokWcGEbGvmuq+AV+88pLPt
KoWPEFRzthY8RW3C/in5Jm0ArZt4C9brE65cvvelXqEsa5cPZkRhufmAKqaYLjoadMW/68FbB5cR
AQC4VCTl2t1ynXLzDAG72djxg2BWNU2FHv3VbUjqOO4E1odC8dlTCDdHhWTtSp0x4b/sarI7wN5C
0j3APSoq8ezQU9M8izS7N3NhyCGJuOCDo89fF67LyATxvdgmd6tv4v+ASYLmekBFcmwrCxuRPQfB
1SjpVYhfz+gpVm9TZ7TsDrAvycCdWAjpnI5QMKNMjCoaDVNPpBaK4jRhE72et7/DC6UtPqVznV4w
W92F6ucl+6uBELhKQ8UhAksRawX38a21XhDIAfSURRonjv6gHIsu8c7PUt1KTJmcACAp8QZUCKtX
3CmFN8zs5/KZ9PxGXFcVqGPrYpXryibG5xtFMeBewN/smbjWQyLqFQEBqjcEakPF4bFqoJbbfBq1
qTgZNny7QFpGeaKB0DQ9BzyhUqJaQv5hy4+LYCfGU2vg50Iavmk73vzjYfEYjf6QLfE9neYxUl4i
hjaYFNEqNKah87gBWNrCE6G+VSc6zHeQ8ryEVPXlNo105M+CEdQ0bJdLCxE5tEjwr8tNDpHL7Xh6
q7u8/PVoF9XpqOlRi+wKKJtF2wtdDqB/ClwiVOPDD6UV2mrMwjeNtJ/YDurO+mHQo4NDiv5ICZdJ
t7Y/79huYxfW5XL/zShViX0+zHI17sfZwzHaOv/v+x/ludmKtYSEfxdmT9Dr1/uJElga6Q11RqU0
HYLg8o9Szvx4gljDC8dx0tovXnXLQPFs8Ge5wttwYhOlFPNMoFzCEfkra8sA/CxdM5sysBrp1jRI
MNR4Z+A3jXQMKH8CAIFunIuHLaz3OcplQ0OPGGq4AzKyIHxcQyBizHjzkGLME9FytC+6WEteOs+P
K4T2LRjltsZLW3xfgJMVLYDmNjUswFd4TvtBPMCuxom9e/iwvaqIktm7IR5mqFfZcMBXdzDZMdcf
n30lEGLdCw+W7cS3x9S8J6oMBZR8rF99V1PmWNapk/L13UoH/HmwBqrpL51OOk2ozSSs+bHi2wvE
zd50luofsp+R2xf9mVBTOxfR5xq3S6oxjc726REwTvOh1Rtv7lTktW+FAkz3hADoKfFOJN+x5PMp
j707fz6ETa/G6T8C39RVysimLO5GZvv3g20srmva6mwUm+bkQXe2bNQmDFUSW/4D9KUealbikEEV
kedYMhgZDIGO1dvQzNl13QB09UiF9ve6s6Qh99xzJkj7zUN7My05DVHo1aplnoqA40YpXrpNxRPM
fmjALMDKadVKcE8GtpaSYx2MWIzFDSXIzMTpH1Ak3mqyif06qqW/m+lyTrIRHoD8JsIcRcAdbiss
hfkttq9xezIWjTBwczLNNKHhtJ+6EeBpbE6BCIPsXmxZrw9HV0cRfp21+IKHAJTDq7k3CB6IiJXR
zSbvp3bZBkdTPdrUb85JOw6hQ1gQK3xS020KJ6IZAvSd0m7firnKfHrBG0CrqIhdS/aYv+KV2twt
A8A0EBgvQs1gRHaF0F3uGYud8kTwaQuct284dnF4bG1SNmOQ6QuYO9ant3nvQ458FsXpoHxFcsmG
Uei7y6OdEKhvxEDFFRTzPvZrIcuDWqKzIPEtEeHZ4kob17FjTpRdNnFkz6Cq0XJvbHI9DXGNxbHt
tkN5zTNzt2owsFzKxJx5qafDRdyrsigAPuLrkZgD/Ucxxph31cF++msHBhwE6qbSLZH8WUiotZ64
e/xcczDVlOuheNqac81fKvcZOqGKD43jUODd3uPN5frgzwsHmIv4d0SyA48kxOh86Ts/1zUME8/z
gVFJDTHhUMfxsDIcVet2YaDmgBLmOaoXZIEFt1GauzLwzYDy9R6rBpLPq6cQpYROmEbUFoGPOSI1
AmfGKJSB+DJOn8xRhd2bv2sAXzezBgjBskZcn66ZB1ObAhHX/qGtxU1xV3vRGmx+78L7yjuSyiR1
EY56Rf6RLiuwKFrQAdWfHmcUL8vByYEjK16pkMa4DaPN3olcERO0eSPsBRWhvEn5hh7+TX3y1WS8
FmtYrnkmH1ydPf6cNW9jpufGN1EgYh0y1GHT8aDPMJXgdbD/sdA9PEr5uBt8xadK6sbsomekIrEf
jPvR16wN9uL6pGr97oJoyra/43LCfxy1F3quL75kjfk3CnEOIpKxetXNKNxC8iI97e34IUhezRt/
ussap5RvmUlSLZyVF2MsIwe4gWA3GD3vIgxhNftOGx3WTeXQlrU/SVVzQ/WhUuG2mgwp+8mrwBqt
04I0Wd4YRpLsM6YvFWqzajnopbGBpr42TOEcvdimYdP6YNxUQaylfAbgDlosvcTuoEYwsTxPAJNI
KFTY8lXmVdY14XPNlgCQY9k4FY4ONdhiAJ/krGR0dOnPJBdvgfhs4qhfyNpmIFECrB6/wdkNkHeF
ln291oV9D/JOra2mco3Oe+dqGJoqO+A8nXhgOpW8KPZTiMpjr/fOaiRuaoNu6UBKzNjlQblwTyQ+
NcH+7vHKBxSwfgxYRLvMLI7W+Kwwpo4p62FfD1Y1dm9tSGdK+mhgJMOSzB5skOptIMyywWsDeocH
qJO0K47uP5tBY4har2bU2NR5vfjYPE41Z4NMegRwMkJkFC/jRZ8pBkTV2gjjWKUnJwtba3asOdja
YxMugjfilRczaIJ1DNQ8fwceZeu7OaC9071bH11yjjKQX/9NyHT9zLGeXFCwQBBGkxUoMeifBKPZ
Q8KCHpH6F+RoJ8SC439XRcU7u2vaEvNnQuYZKM+R4O3oTmvw0mG49ZweRdVwO3Qc3nNfUWPW6XDG
cXhat3RvA4l4j5R31SedopWyHr60TuMEJ3yZN3/0rOQVdS0gAkVWThP4gg++QczVy6oXZuYzJaHP
okTeP5/ZgQTLQc56tHJ/3UKduRbT0NCV5gtdAQVoGal1U0sPstXmigDFsYMvcC+GayYAaol7V4Dx
XbiC7c6ky8oIayGxb2AaJwzVs/5FPKe5BlmuAp1XIJwfNtwak6fCvZlXQekZvXKfkqeI45rLcQTJ
YB5Zur0YYmFLw17Msoy6wQreluM7VFUwoNte2HlSLbC3dIbrCrUGLw8w3RPQofncj25a4z+K/9tu
5pFUEWHeL6Lou1x2JiCIg/g+fEScIS3mPLlqD+dtuRhScTlIK9sMl8gV02u6gN/iACiB4+nBFfXD
8L5nUnyv1Znhh7RB+M0jjUfMHAy1mo7xS8C+udXslHJAARCB+tKSAjlxKjrV+/Vxo9hK5urC324g
lA42efYDiyq+R9wGCD1QR2OPXQGwYotsn2CL7LpGmhsZIbfzmM8jyYloATYH9pf8elSDYBADr8xN
qAK1o7AoxWAByZJB3LG0AYxY7sNo54m1yqs3k+LWG+lyqPJhz9Jnupn/1IM5qyagr0xfBRC6Lfk5
Hi1aEo6fU8FoWBQ6KBY4YPHMHmpgz+wFCXmHuVJK+nIsQFW1xv2sm0Xrd+5YtlV4e3DgasCB2Ijm
xtFacYFoNp5+hQtdONhC/K7LddFfdsIfa+kPWiZlA3IjU+QEf+QSrUxIjEzDc5Px0k3sr3DYY4dV
tdX1jzvNIx+1sqY8W4yB3y8XXOZRhrTeWAomS9z7O8EPL21/xxPdh6K9sL4e6r8hRkdZvtdF33NR
6MJ/cjlNBXq4Ndl+05kF8mxgo5yZWVN5c0E+B/s8wp5j5AOpFpg34hXMVMKLuuI707NBW+S9Rkki
zGRZ5cX/aRs6FVg6+uAXMPaZ5RKuJAVECE6886XIsNSDye6EP5W3T52yNA66R5B5u3k3uToVTxK9
AMvur/pMNgfogauUlcyk/QcXQvXvrlLIQr2sRAiR0L4va9Ux4Er8MTwuf8U7AmB39X/v4duOLMMZ
8q4ZaPC3QxXawHJZCxsIkpjiu0gaZbLY5s8bDTODRDlRzTZlBo6oWt0PkHcoCZkpXmnhyNkPiAVt
KY23AcVyv33m5TN8wk6OPM/w/JgmQdodfQNtWnrUkWyTbfhV+grWObDqk/ZmXwltHv6VzkCiOF2a
XOogKJsDIsWCgKBPVHFpaEgIx/3UOyM/9ota
`protect end_protected
