// (C) 2001-2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
mivzB2v23vktPCJvjAr/Bl5V2+CcDOqchiK9u2xPFXIU/uroOjjVZEq73sRiQ+dkGUkv5yo3M3iC
cOIKcchIYJNrO+G5dGzb8e2S3zkt14/a6L7HsFOmyqZEZ1JioeGZDd0IozNurdy5lnP8AyepPpG3
O4KvtFyCrfkLfShuscv/wRhobcSMCuupsfXkhBrBL0xWX4OP4bvqe3tJCIpoL0I1VNnQn/gS1eaT
u6IBYRDyaDP8dKdpc8pSvIN4bmtedj3yK8SS7TIQvNZycKMb/GVhPNgH/lMoJwiAmOqDCI+aRsD8
jCEapm+rNATwf0znKRBFWbWiOWTyOOFY2RAiiQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 21216)
BvCUjQCSdV3eCuFuihjPmXcbYCw1vFTUfHOg/tXHI2LZqi3aBZ43e4eqG8vhVuKgURk/ggrlU008
TI6bdd5O/vQ8O3Vi7ljsL80Qpzcv4RBe67ShWw61feMKH9+/PBl2t8PRXfwcp+EQOF22WuYCUXsU
aU+ohguSlbYaTuCmi6IGsiZAJS7vDDpCfS7qKrUt6aVzNARAlrpWruLll8Wd+jcEtlrhFAacXYdS
NKjYIuI32clSQlBW3AibH5+BslvVfEZAZDdJNKqC+k/zs97zIw7cVCfERfBM6W7WMqffPiEYLKLk
1rWSIMNO8JA/lm86Y9roATYAdyhsEKH2zH6REdLXI3N9f8cMA8XwAGJwWGztxi6BJxmVuZWYLNog
gO46QzXvtrO7S0QSjHDYP38hWosAfAFJWQUBuuOwcLLczqWk/qzCZL7M0qLb34TtVRrwTswIDW++
kaTmZUa2LP3ZgX25wAVIYpvS+BMgl5QXnsrUUc7q2ggjITrrCYVgpaTI/8lFlqViOUb5UBVvTTtq
Zy6yfe6ZEx59ogQTmVVEiy6AC+B2HRWbyBoCDTAp34/JpDwTNFKeQX/uPBxI9Wijwes0Tc7eSdvw
/92eooeI9k4vTljSyLZGETyHTeK2YXLosSeKBxtaW/j/oS1tk5MS+B3drIU9xqRL7y8qkMSF5w+g
7Pf4d61+NAdpaT+IpfKRtb/xC3t29knHI3KeIvQqaChJXnTlmNWXf+wvzeR8Q0JfcUJtOe8JbYA4
iqqbz8fRiPtgc0QRT1tcYAGFUzEQS+YcQOdefKTUx64Ct3fzbfJ236evQSKVPQEOpa6h4v3+JwRo
JnfdlvmZ0bHzdjw7tlJNnXfeLDbk+A9p8CKrM0Lt1p+cyF/1FjcDkYxqonV+Hni6fcxRV8Zlc/4D
bq0R3W5EckA5zeQBW3dCYZTlknUTFjE2NpLQoEIEDbNIka0mvpoxMLJi/DKaIPigxJEV43WqGMRT
LsUJEv4GzGfqicOlypuad8VG4GAX8vypI4WE2ETbrwxwLzwUAG7GFSGlhbnlJbRzjvoXOXC1LGEY
R2WPTT9oakczBKx2jZG3o3oYzjjbRI12ZJyi9jQMK/7zaHMikGk1pkQ1203Z+PhQGiLcPxsjjo/k
6CM3r/dLOuO/yfii/8toGkl60pveXCslN7mtUeuMcNxA5axVD4Y+7Q+cuQKyHi4SjCahCyS2RBH6
Flgv+n9k++yPJuj96txK3yhxUJ5VRYg2T3mPGAKKiMRj4t5ewXFuoCeV4vcSi5TJ0OsrCvDV1ZtP
CCt6otFuCRswiNjcaIvtRSpjJwUYfRP5NPmtngnGbrRn42Q5J8UcwcTYqUdt95tiVgZXLICbv7bB
TQ2pQxiCXKJIxwo9gMlysyP1e7wNP94NmT3FWW3wKQh0QcvOZXKhQok4KYBv7/sgQZ5gBRQGY7U5
05v+3HPh6/qXPO9jVgUG12/fWynOTX9kOpeMuNvLUTpkzgtlvfwQfkicDQE/dLinAMo66YKRugAP
s5W4xdeh9I95AAoxMMHhAjCNCMCehGUNjVa+30mGX+YDMCYC1o7XxFWc/m1hdgnl+417gkOK7lh8
3MyWLBuxG83SmwUijFG/0Z7WGIA+/NkdeHCUEVN5Bk4NurEG4nZBLLXv3RgS8JbtnWvd2Zzkz3Sk
Uj4zsFtHZWSCiwm/sMGfqjbQiMWTfUPr8V0H2eLH9Hg9LyoAPP71yLO7B4VM+3z+LU+TOmUkMo3j
rjC5fA+GUGk0kJKeKFg7ldq+AaAoNT7HEPVL/4dARVgHo0T91PS16kRNh1wjtIavzAM+pCX5dJEs
iRUUEOkjuFxqtbyETrgHcxCPG26HC9uukSn9+Z8tZ4DPELnh6b2gy9DqqBqFD/eReksX5hNdY3fb
XkSnmku9QlP2jixXKI/nfEG8VWUeuTutmT2i9LQPVHV4B0DxnNGBXODDmplag5bB+Yk1rqgifjwb
mZbnzrt1Yo3z20ybE/aXaria6bMilL32fbcWoKadxpx9HL/xPbTzdgbq5RJslJ8IUCmuVnwjCUiG
iWk0TfmglGhFpGY1++uBeiNbLXEvRH0yOUrOW71OqVQwqyooU+GyZpDmZqozBMEPNZkMLBPMw/26
sJEdQGqIAHBFHpsFaWV1l1/J7AF590ccbshRBDTHvyMFuHAy1DqVSvejFhMF3IBDy1DEr1//cSFM
krlkjqmB6ywyY4p1HdSsNo3yzqwG4svvq297QTLfvH6oUl1asut2+lFTqkvpjMJ8LyrrpXR5w37q
Q1fvaDcZyUNLAAwe79YCUnHkGeyaYq56O1ZNV5G/yLsKrzI2R5RHxXpIVXpdCbaAhaNLSN5XfQw7
rWGoCi1cV69S8e9ufbMQIkvLmV6rRWFnJVDqsP26GV+IVkrlb+tMEEOlJUfNqUgWXnwfJkT1UoG3
XMbOOQnMhO0PMOGccLqZhpmXw/Oh3t2qxhyvotjCGXRVOjZlkKyjM5ZXwzi6MHp2NHnkYABcd1AN
CHRlim3POuVVIds3bzKRP22cH+joH5aSm4fJFjTUXohspP4FxngkFDAV0Qkn4d7KHvosr2I1/EwT
5IfEM6hjMPyOv9j3Ae/gC8+FqM7B8MG0W3bxHnnKJVh6/CfxCFOb52jHk37LdeoVJvZXK2xpUN7H
EhFgcg5HcdYlO8QPup7bSrO7u8Lz4AgQrE3GywWjIae0N85k/PwWrR6NI9RZsTCs4LJyexE1CKSF
grjiK6rrDkTeY3zZboDP8gqDppjLtvNo9NFkncTiPMx/pm6RJYLOMEHx8WoUJcYchzGIqZYe2olC
wgqnVlQfMURJmcVJZ987glw/AMzBdGeNmVegOnQBJEn8Ug0T5eVBue0ORiPNJYK4ZWyWZm4MeecM
eFvLlksRs9cqt0g5m/tuRqId6KwavgKro9VzLRh+EKXdO45GDxwVDtQKp+pgz/5yDJ4aYVbWg/KE
35HVbrMg8NCTlTfIG2Z+Kl0TpDBAGAHE822iO1NzU0oDmoMDOXDl4sS7+IY9x0Ppvpyj06zbvctA
2mBNdd3gXnwn16sYJY5xGFBqHUtqQjSErxJJVHKGy3Z+wphGVlLo86juzaWb+8baGTOVXQBHB7wd
PdaqhQQ/ejvBp2a5DIxN1nh2AfBceNlhHVhzqz3TSSd45M7tYKuQCvNy5gHpdNjgie1VQk3uUtG1
0eXOEeb20WxuJ0bHUuIsNh7kUDhQuoLYZHnW763TcTfnJ0PU0ayc/cxSMRmkX9VwL6LBptwgSajQ
32LG2TglDlAUFk62en59O9k9WuTHaNouq1MU2LYCf/zZ3m+WgWSUvOKVkMziHziqII4tIGZRlRHR
Biyomo/YbauT5ipFZ3SsK4B8BDgNA+eUDVlByvxhIol60sdAevkElD/HOdtSpKxsJ1v6a1OVJsFW
I46lIkh6bF/Bs+gHufsWMPgdP9YWaV+R+mRdfZhII2T2BsCKZiiK5o5I2nRRANQc9lek34RqIbJZ
quZcyLOVbja4y11J9bO+fpguW0150XMGjD/49G7nKuN7VL2GHybRDVHFu3v9ysgK/lJFrmJwwp6o
2GfDgpyVYZuNoHgDn/u8hqIXyM0HS1LoaZYoSoRtuV1Bqk9sw2jUy0R9JiJ0tJ8h3KYEMksKXj7E
ijN4WemM2l26cYt3/PcLhcuYwqTFHzRoKhKK9RbnyjninosfuT0KLByBuigdUUTza1eWFcXTOAXr
bv8T0OvgdyTz8nRfYggNIYpi1RnGd3W/63DPWmFA0+RPd0G+vJi0cq/QWyotPAOSVj0jLKK+smBI
rYWB8tutj7DUh7/4g+t2GhqB6WGGWEhiQAIJMPmwqSmv733g0DEf2bS2V2s6N4iRQxmRbyLAtTLR
mnwWpJq8Ba58GxKgsaDGqBLeacdnCWg9ESd320uwTeNFfdwZA0U9G8NcMPYZvSZ8x62XEiRjLDHZ
y2PiZ8BueLQA2nvKlteM0t0oHtF92w5f0fCuftECjDJuIzW5guwpzcPPgz2HVkpS0atQJHMJ5xSC
oVMuc7KY5/U1LeVyNZor+MeBwLEAS7jZ48MCo7RtElz/c+RW0WujwRC+Qbw5/MgdzRyuJRPUjTtH
+XcXtVKhiDROz3cj4n4LkHwNi6zeSjJ7ByNMSDZuAYudThazyW7dXwWPHGYNwEJEqyG4/eu/s/8k
tA31XBVIZhu/VHDB2qMv0DQOkp/iIAfwSW6LCBHKj/Mu5YJEhPvbP924bdLQksPPYtQc7iEkwMsz
jULmjxXFpPGf89TtJTwu7cZ2m84e5hPTAuGM+eP1/ftW2v4GfETB6CiztkMGZCr1ONCYdxh1broo
eXN8eq/b3JUnPJuVpnK+/2xFT+nYKmafDs9V4cob06SXRrAkxV+5aBhp9Y0HZuxzsM3WLKua8Sq8
QnYCGTB9iaZO1sB/9ALTvC9DaoxH08Iv73IfL+DYYIyQRz6GIoo+UD/Xm4tfs0Qfysp+eKFADGjc
q4J6lkEvqrDoO+vOKxag6NN/DpluMvxhknJpyr+sBPauJgqzfQBmx3xzEc78XqVb3NE5DkWKCLkg
BYxPfHsMFuWMukQRgq/tVEeUcYVy2VplaEmNteXO+2jVYsjix12hjB6HrhVAWP+ssedcyNEBxIpo
UUYMCwjuiW8vdTIe9iesnXXwsq9vSpTjfzVL1q6k92MY3U1Sy9kRB1FJawBrJnYsGzD3wtHBHZFm
HJt1OjaG6ELHJJ07b4/Ze0cyxZT83Ve3TdR7Ssk1w4sZ6CaIDMt/4uwc8zxf+j90pNCEOfyNEcgb
E3gOx7OnxIzPze93MhU4Sbzjr4e8bHWQABPALH6Gqp5LQJj7899Uyyb2xz6FOzUYKAfk4mUvDSZA
1WYe7u2KC98FIyOgCwRYntxtdkNtO2YYcC9ZMPIlgzQkAH9QRghdqYGpbGFj+FD4Sw96ceNgjiNr
nEFO8wzk1wSspWYPQh1ZzXt6Qe8nT0A7kVtWHwqKqzy9DaM5IWc7YdktClVY/s+FKzL7BWc8FVuX
FuV6eJLEjH+SviyS6c0eBvAP0PegTacFOBWyzDyG9+ByBsxi0xPemW7xj7ctYiEZd6z5+34cBkRc
hLKkZ6HirqeEDtxL+LaE4+REXutLyFa/pwlmP4qX9Dp0upgsOMu9CNfSb5ZZgT9LRXIHyXHRutkk
i4BZQwnsjM6sXc8eKGRpCrDe98J4XK2REY8okWC/LQFE+d2VGBFII++36/ZIdQkb6WApChe4iv9R
Nx9HClT6MlzWVT9YEKFecdSQzYb7vG+BfFfK3u+H7mxRisv697s3DY62lv1uf3BOGgR95LG7DRQG
pa8RXyHpJZKACNjs4OGzjvLL2ZG35rIaPto9isvFXp0Mt4oKeLmyPYlxlCtIHktQBxC1w06AEo+1
pENBp/LUtO/6nMPt1uqoSe7vH6iM9JXE6g60qkTwTnwoI0rAO5Db9qkTirhjkRjUXYBYrgDI+FhQ
DC0TI/QW1VwXYLjIEY+u973mJMBDcf70Xiv/TJS3lYWarfsMkvNorb0c4YCrqSIu5irrD2bMydL2
Hsw6nRb2ftmk3sU3RFk/eSWu5QxmL3REZV0WvifQFsj0ZYkt4pDlm7MNfe8BDKGTsptmNPICUyhy
ROBw2fdECKA9vHkBgxPfPof32RClKf06rCJ+QBw3rhSfcU/Rr8OWVURB6OIsXDtJ6U9+xdikSGH+
VW9KekzbPIV+Yy1Z3ljZoZQgtcoVVIzskOp7IRnid44xhScdLZJk8NN7eVcrTY85b2P+0YaT6g6W
pujMHkuHPk5f5F7whVfYkf0MlL/PYzs0tWMg7kvJmuvXnzT8renQVJvi3OqCFu7niJS4b+dQNssv
Xzub0dzzP98Z/f17fbTbn4he4SwVDrj42U6Mamnsq5WOxDuGrvS+wDgyrRaX0WA+8Snp3/MAto9d
1ox64lA2/WCw03u9X2nrXe2UeI0zUg0lncH/w0SnydmVvvsXrz/+k6+uPvdYoFXKOQg6AZ73TevT
KGMC9xf7CB28sDxepbuyPCUqREo9kYyayCnNgR0/pyV73mxxhhnlsOGR0yZMi0qbrQgqasBNpFf7
WWLrfOEa0W03Zn/gPwI5vcbDDrZB8RtgNNXjsHq21QEqxZAtfXsnZU02eR7vpdQcoKZhb+ibwApM
GMrbjI8KOUlBVj08BU22YikHlPst2/jAtKDvsFJiITUH8DM1rWx6vfYaJapLR1WAR3AWIHiszZKC
nBskKlaldBc4PX2FEmqWOAbkBst8BQWnWf+FgqREcXwa4WzZLtyU0pJKN6ZenMUNc8eSCTIA7W81
S6CSzIn5KlU591NF0FB02CpRxekSwA6mWfFEodBZK4MGB0VJZ8Ndf8iCa1tvl9mDGbF9aP5Y2v8d
gmdD9iZGahY1UG+FmKM7xYEeskfExEL8uL8dqKvmhehgND2joOWSDt+li/CJo+CFUdEDDkaMNEyO
bdyYbGL77UIuzDMDWZjYvfu6hvtjsqjba+Fvc8Ghi2WNO0XUekIopr/XXjzcJmT7YegKylhFIkGt
QMU9NvQm649PQ1LuPcPEkCUrfhDxZ+UoGWnoP4+WhjCBlOK+2hpWswK+9Il22FSbvPNZEb5qH+dR
TblcFQkGTgfp4QTlH+SYP2bKiPVg4CE0n2HoMarOlTpaczWQIa9Me5srd7dyBf3wipK7sCaCxUuu
g4j7ewbgYvVAfaTs+p3jCx7mfkCmYmgBbIBqAjWx0Iq7Q5JSZiPcAFnL5yZ3MWnPeXeoAbfnLPW9
6L1ssvtfsqYDRal+rRLazoZLcsCekhtitBcmuE5I2rAnCOdYDsotYVRjWmLMvP3fy0K5ykSK6kQn
CEE5yqCvEB82PArZQWMRYoVWOKrhWY2K113Tr6Bu95dFuhPnI6BK/M+QgwW5jdmzSZn3oLzpB02E
+p+dYOj8j15hImQXQKrk+IDHsyD4pb+WbKHDJFEZgjt7JVbeFyrNLTOupevyh6YfRWodq4jHeEua
zZxvmKK+0821lpfCxmmW8wgtbYDUxjw+vaxWFl4jMUs1QxRgCbuRYeAdFMaVTz94LLFdq44uBJUk
CSw9zp+wvmW+7T/Mf56axRMvm9ZxZRksehtV7qHTogOei4fhO7VCRJwJteaVt+Rw2uJV9Lcyz1+E
j1LgwuoXBZPN0ebmjEfv4sOo48+iiUWNXbPlN8SqyK4QCCO6Dj97LqzjTeZ1F4BrvaGkfytTDoau
Pe5xLXmKwuvVgKaVW3jEW16FchYD2X56uireUHhhI4VBSA2NQGUuOq7cM6ElQU1QdFc3pWsTXSlH
kMy6EiFCYJkwkAUHqtfo1inusUCBrMiPfYvKGvbl8zFqDrJ+It0jEnHEaVlmnqYDQh+vOANAN5al
Wq1PtLgjwOVa4/vzrrBzBbJTdAr+qstDhmUiOGgfccoG/ykBOrzWK0+BWBH23BEof39drfBB/pHB
EVnIIbKjyNp1LSYjnlirnZ10VpG390Uzgj2YnZF5y+dET76b73sH/yZkrL49wVDqVHE4pgx18QjJ
qkLHKyZWSSAx3t0J0ToakieAhbxNBTykInXziZlisPPXALiqLTywshho9JecnNT9azkk3BQwcsbO
zUV4Wv1DQA/xDrx0LgfVwKmZcX64fo2aO7JC1vlszLF+0S6Vietfzdsjr7+cP3PKiTxzcQFSBoU7
FA1ZNNC+1EvgTTRequxBO/zechaIg+8SSlZ4SKycAh5U1kLqPdylNBkKK1jOvHV+fcZtkXAzs7OC
9ggVndQlttrMCZI3nWKq145UaTeU/BXR1FwpMUHRch+gbz5yjbmSblD6oOUW6dcLCilzCRQDGC1C
Hq81vq7q+IaCRAPDoWKTsL27wB7uyrTJqshVhN1gHKNhxZeqPvRpfousMzqd22yhMb3BsQcWe7Kv
Ok9TR4E35I3ypwlnuvxY9qCvPdw/boMeEA8fRDt01YIQXwXXe1nXgIMlJE5w4AVWSEQGB90NXWg6
VM007qNRAn29aLc1uPwjAWgasl6SNvuZJbgcSjpdBrcrBw0h//8rvTrUbuIDlJDe4M0/r9cayTfV
EQ/B6gFfutYA4e83ZVdsDbIODiW+P/AvYLfzWRfvPK/WlMAj5z1DB+f2ZCJZ2Zh4kwLqxBPWQAc9
+2gBZaPOYlZ+xGSNNFAWe1cYP6B1FQwksw/hGuskafeAJEg4sTxoPh3UukfCjj0pv1aQiDKlpOh6
8MdiD6rT5RTsFzihOeWmbME+Swk63YAeuApK0W6jdR/Qrt1yU9Gp+LrxI/gCie9eL8CFlz2xaztm
Ni2UCEP3usi0fIuH19SDuTfUUKPjFbGYuOxgQpZNfjXMyc/7nF7wFmNlBJoIIahEd+Xy1p0N89P+
7Jj7O7o6+FcMOpnqwYx6GB/s6GtnR+7dlTs0czZbpw9m5I187RTDDdHkySqkhuiyR1HlJh0zaY1T
Ex6lEo+1+bRKwDIqdKrLk52K+eqt1ebS/gZnAPBWBu4/zDnx7jmJ1BUAW6518zQrhq+eq4bE/7al
FuBj8Y2PbJOtvsKDMqqcTwi0GXbX4dMk41STs/BFK6SGNW3aSovCnyDNDgj/pSw8lJ1/Bcrpi3oa
zStD1SDTZZf4Sjf1zqbgHSjPejY3dHP/jHK6c76YLJx+yaamk5uXJLpBJWWfefUakj3sVqoJjYzz
xrO3ZoEEgSq6CiRcoC4e/40RzQ02JmBt1epHailg6xtg1kJfvnH+DI98e0OVc2sl5PY4/9b8DTdX
gKrCVhH+R8ikwDr4Ok6PAsSA6gr+yv1TBay5fRgIUPww05xyUKx+9C1T7wL2q18lbbcpiPSzE5r3
c2ksujkodFLn1LCZhimoaEByC/ppsFyMNMzM/Dc3gdxC0Sdmwq/ZQ1rRwzfL8ZoJtzKHYR7vH+Vd
eXhKcl1A4HwWswIIvARX1i2LvCdUFNaPVrTir0/zEP5Wvdw4bcbuU9RSyGng6NvcThf6rHtarveQ
8+1k6zHOetsg/ijsgm5lIYoHYuU/cimKOFtiYaGfdhy5zype7z36bwork5T8SeFUVO9mJrlgo30h
gQV3UyvfCF9TdfG/Yvo2zZEoicVht5ZhdqlqnVxHB7T1l9GE/eB3JKjFWGvQfbGM/Tkka0Uhk6sa
NRwo/IHmbTLyPuVUkwJuz+R0Ttq4vylO1GNat7TyGAR2bPD/3Trloz22jS7JR+jsPgE+ROFlu9by
DBBBmXNIJbhC6WwZXZwQmESj2ccJFPaZdkN4qkSYjiVAjN3qSKaQZcJQhNXH29aBSSoouYbkMu7f
ygmc0mVVrPMMzaC6IgTFbYQ/64F0p2rncFgQpOOoePSqEEP9ZJrTsbjYC9Cnnh0pOdVfFOZCgB6g
v6AyIXwJR6QOhY59W77SL4pQOLobW08EpjqgCmZmDAA2lisBJ+q+J3Qrj98uKnqlFpUWhkgJMu94
I5rkr23JuNuhN9X1gjbW5VYu396XVdDdq5k7OVd0KA3wm+lHXsfFNoo7HpY4AuFmGB4W2zz97crp
zsSa57AoeiT1+3+2Mj4v11REkbLUjbBxrMCsMwT94169swEv9N/FVpJontm2wW+FXZYxvg8AvtkG
cLTV+mPHJfCnpCHjA3jBKsKY7lttiQ339/mINcjYsKWqbYqhSKYqc5eMxYw0c1ELi0+CFD5VBgAt
QXMqA6c1g9zHMrYoIZl4819s7lOQgN0d0izLrpqpgpsFdXzkDXhcnyGl7a0DMsDhPNTg9sZ0vwAy
eajwKmOyyxwTAo2CQ0XHdliqe/A49L4B3DlIu6XjcblWlV2HcD4mP/3QxWdp/lJicvRPbcTm+sor
c9SX+1FD3u9yjbLvHCWcUDW0zHTZPr7gOt+BdgEzruDZYJUzWIsXWDswbclsCu5wQojcr/7at8KP
YxRle9M5rPXD5xQshQ0lhgUwXOKasztPXZ6pICiAYkF9L1FlTVQVANjNJOspdNdP6EfwR1S6hoTg
0LR4f/jcv6cBSMD17mDo+2N2d5w0tPYaGdYxGm247x0rUwg7xQgwUjrGjR01pcBkrvqkD6LQmH2+
9IViLHaJ5vyb7k/19dOT3fEO8ERqttXWcmxxEtlpIGCO1Z/igZvJlDjsTd4qWiwJUoh/tqWwEEe+
GOUk6VhZTP/UhoUeXspQGHSgnOTiqGuE0Dm8lBu6cTFIujkOIyJnmeHMv2ghYkLw7b7N4F20WGWR
b6ymKqOrPhocwq11X7pn2ppviNpHAJc+0F9fPzycSDwS1NGPLswCjL1P9uaU1W75zmV1wPemliTS
jXwPda15W2f71CZrxQoZBb5oj1gFfOB5WUw6tTiPOUNHPCNB2BD3FXlZtQq8Y+guqYyOYCLiTn6n
jDBYF39IVZMJ6ZZdAoY1stTQZ7lIz88WrWuDwhBESXOktJf5FkMB8m7yeWVsRrDWwkz/HYEbFFt7
duktXrmTFQkAFcGPxeeq1C7C+nqJTtSqDgTZhE8+Je6ncqK6hZha11raNwUGGaoU5yvXYmYtkMwg
hmnkPFIS5ti5aGlmS3xUtEFE18d4awU6I6nf81d4tiFMsilhko4aVUvfnEnMp4irxQP2+9v6kYP1
JcCaXN9csAV7pNfAYTngfW8ugn+obMV1NgDFyAbHTe5EX8MQJ4jWJM1y/nJZInsEO6aZdN7H+EfW
uU4yNOZSPbO/WwXA3ZfYz3HcK6wpAqN7vGESNOCn143pa3sPbRYQgpUrBvXkxk1fDXUYXmdV2/0F
JQ6wSN2GXrlGl+efWQ1eNC7Q/ziO75nf9NpITgcdrVnG1NscQ2KF1ZhTT55O6iwB8/C7A86mYrCz
jwNFb60W+Sa6+oAg+xnFPZ2dbK0SyPRczm7mGAVqAirllZ2Sxfvlzb4Cki2/BqnmVm05oE0iZQoo
/HWYI63i/TQjTBk4afKWsS+BzKY3zMseJdu1tnfXOXhoPCHjAb21xN99npq6XgNzLmojfNDj+u50
EosNJ5eiZJ9Fke/+hDhALtPZryWUtCZtPfcCssAwX7G4r4VUDBDMJ6Cbhpklqdp2WhwmOi0DEqkJ
K2xfMWuR+QZsl9SyNlmQzgrCL7juTMwk3vzwIU205jLCDbBWysSMed6Lz+Ca8YGoex9vPPNtH+xX
pdb1qsItF8kBI3w7sXi4c6BfVCdb7ziSErF13FvAcKaJLrHhbf4uP0JMA80681lOyOTVaOTxI3U3
KkR8r9l04rvRTQPVsvUVQVuTJQgeXB1rfGrLswrASv9ZM0ALZ7ew29795Wg8CZuoItCwncd68JVb
wIsJYKgZx6IX7uT0uBOZ/sKBsyHb7jUGGjgtcos4L+zDrh8xjNDqAUZyJRXrgLqAwCYm2p3leAhQ
c7YpqEqMhZGYrAOajQYI72zL3DvQZaNFNuTAwcfo4Vqx73l0HnuX/NN34qJY7tezBI77I7ZIrHTq
9Bpdo6MzxVm9LNsBEYYO6w+/SgG86XvqrqTKsgKD9/mbUT4KZWL99sfTtC5A7k4TeQKWRr1Ud6yL
WY4Pzxtp+Itl4FL3m5CCZoyO16Ksc1YLQHTJaEEFSMA1XgKxKtfFSnj+qRnns2hja4jixvU6scFM
2dH253j4tU037RKwZTZl2pVMY1AVg42bBvHIuUnlhcqUp/n5araWjLtfsBkBvs9UVEvW0EQsBoXD
kmElifJk63BR3b4bkNqI72ivNZW1qpUse/wbcjwDK56YcSXHxVrbxDnS/QuKjfDLtudK7XaEYBEQ
SOG1NCetvD6cTrcOarlU4VlSkPlxGRMrsCaoFOAfLf76TpDCpaRrbJEw2Jeg7tqNDzlOVxv1y/mD
99UbgKO7tiJabOQaiJtU7pepvX7LtV+ZvUfAIbZrRSXOA8Mo10IBnL8eQrgeih7tdVMI3mq6Mq+w
aoD2mgZ0beaSRcwGG9NhYCC3x1Il6FTCetLNcalJMJhJKN/7LXbjX1E/hDDtXd2xxfre79kft4xu
T8asdJV15R+bkQJILcf8jYyc/sN5pTP8Qjr6TU7GRhDEtIq9LfG+vXGx69gURtRaWZu/T7Za+PQf
7QA3f24QfyjZPBO1d0HNWGsPhOwyRY4UPnTXZoOXt6nwJXtcVCgpSdrHuXqdklU3cTwtFs+J0Q8i
scogPlTpjTONzpnqOcv4YDlO7y/4Vf2OP3B19f3MtuHsKydChlfUk+fUbaiblQ4k36bhMMQcTjVt
299mDI6bK+oDF1CYxgBemIvp1voAIgm8tIGv0EQ23CZFXUGpXkqbfcAjq4xHG0VaPrkxPdBLBk/j
SQs1JBg31H0SzMk8nxtEt+9UFYentWsFvKoxmKTgbxuajToV831gyQw+uoOED85h2ebm6uDXg+S+
h3DaWDXtfUnmjXDu3xGYt+AWFf78KWxE6X/B0ir7bTl9nLvO80J3col844IU6MsCJB+T+psz5jTa
3zv5AO43hKOf6F3Jw7pibxAN460z/2MU49cgYfTgjuhSCMFUiB+CL/IFOQ7se42G4yX2bjaVKMAE
j1NZ7Yu2O2mqWO5C/TmcvezwR3pfpAdz9lKB9/N8FPgIAsBhjGATTeRVzycoPg3PSqk1kWYYoMTR
SgobepcsOPEgG9fE2eDCMBQRPZFExIboCtmWSfk72Q6OcY6qdWcs9nsNkBUdLUVMPsFTQIF7KvtB
p8KoFyO4HPckEdD+chaUa0vU7U/uPoe7+J7Rk6mgdA4Fq8R9+gherhY0ar4Lvy7xzu3meIg8/jse
GJukvIyQrRxlnyU79h4jHkaW5HFEw+9Pg/Z5G5tkIyWvsX9bmzVY8n79Ct/9CTXZn6S/rfDPvJyT
4AIJx5Fae9qNt0OvrAObT65qKHWoTnVU/TmSCpZoRKIQAUmXhd9QaaQsrTFJfjabuxloF7RluheT
v8uRXBnDIDyEarr9ZwgPrcmAb/gXIo2uCgbtZPuGOb0aEmkhbb3QmPG52Qg2JPdQEaavvM+ZdXyn
W2HIUvn/A8kA9gSLCjqKKgFw9NEaCJKK6CdE110cxn130EgGMTTzE40raGxdcd5tMR4FOchOT2qT
qkjCug4ya+/dIHz2Am5pIiEVnAVwRhqJz5EVwLgIa70ndvV9Tkbhd3UpcvkIeDi/+9W1YIDwYDz2
G+SPPIXtJNwK2vokPKnjse/s1ksT/965WlLcGpVI/4LsbhwZErajzB8zIeMhdvkaVwaOZS954Bfh
7Tgm3nkE1bSy2GcSyHM6yV/vb/JaRg2DA3ThdnHbDDaP6fG0FoZP8bMpLjMX5Rdp1zdZjbr+SquG
anX4hvP6XsXPkV4FiJtyJ39A+w4Tb7DIM8HuWR4UXLB27AXT7BiDU18oWhBj1q/J7QPScrWBiHpN
kCE4dDOee3A+j6Snx9HzKTF/BLB6g81HxvkbIwcrPuiFC6GpP/bZrOahHKP/BfQ8xkQL9PvD92u8
Cj1KnZ3EsnjWuKiMBUGKzo1qe78SIPLLN5U3lVScjU9jpBMP1RvLMoL/Y+ckKWt6G7qpeiWQhSf0
ZLnlBRHtJ0aYRH/yOkgv/fZQXn43uBgVGQIVGR6CkVS5K1AIC/CNg7kWhW7gjTovbOY8AuNiE8q5
uhqh2xRzjUH809lKKbmpQ0HGPdTSAi0JQfE1MfGTSzh2kAYNzyRsmz0lA9HrM4z92Ft2oP+oryYL
Opclcas5+BHKC3VlXK1hY3Tkp9294DahNVUPSdaaCr7WGIPZPthqWq+vwDGSqSgmCQ45Ze4zZzjQ
AQ1xc+KOMAawx5BSs4zDCugW6qRz0IbqgbA71brI61SyPMXHEwc7YcIwPXq6BzP1xlHt/edMihHj
3hjsr3MDNA6K+q7ILnXOGX/FNBO02HeRTYD4LtpHvyPezxVeC744qMe8b2CLbGt3mjML2QvlZ54+
eJb0ZA8mImwOxERkrRmIV52qzw/9cT6/9rB2GDxed/DKrh7Ugm37zXD8zQ1BqT41dDeoT2d+bdhU
uswY3HsdChfn/FDwcUloP71V2cClWlUSx903tyLtjFRLz9w8j8KltV6oTkGNjokEzVLuO7pGid/1
+uKlEjeT3IPF1xnMHWE0dARM9/U+gLV5HUXkHgWzClaaX1/zGzmMk/1Wv+Fu/f0piosrhfLsCrYZ
Gea64kuXXrcvrpyXuVlAnM7/qj5MDEVlQU7ssDIB/WwnkNKlYb4TYgYgE63Kh26IJMqEswKydl0M
enozneGoDk0QFlrBNGcdHdK77GoVE5RAEh2NhXtLguqUovz+HB33H7HcCqLzWBAUeex2mVJBLlsx
zwHL18O4tu0XdZVclo/Oe0VJLU93Y7+41fTJwgWqfBdEQ8o4wibbxzQwOIAtXSF9Y6B3xf4DlrB0
FwdqGqGIo7qKGQbZzjoFbKG4erGtPLbJU+TRjRp6Iz414iYLFSGJuJFgmg2NlXU8LFtk+zkV/iPO
vC+D2NqR1Ko3G/OnshV/dZzcvjEXkHIWqm+XEeiapf/OHAHe+xMG1L6LAumrMum5rSpfWQhKXcaS
39bq1fhCQb1BlbBm3Qp2grZTbhctOeheNb7mESlBua2ev0FXRMR0t0qGKoZYJ0UM9z3rrc+bZ8Ho
oecjVjLpmxI2VEhXvl77fzGAf2N/UJzAHiVeZCL1rhc3CToOVpccBTk71o04P8SYhPv+WEME/m+z
zKwLhCD1CtgT2wA9SaYWDEVzn8WXa0TsBgCg89QOuTQlU+pH2DJQDW4jfBLSs6sdfEvM3f80fZxw
TQXYMABHjcLPrjqs5FkwtO9Vqo1RHQgNtbekuMW7Rh5Zz+8rvrJL06+oBEzg2g5YvKgExolqnFkN
DJFLEUJibRQ6rpKrTDIVXTCdbKuaRc6tR3FpsnPvm2WPU/IeGNdJUDZBK2TZOjwJjT1zM45+OCQ/
wYD6PfdItw5MrQ2XeGLGJoCkUpcqc4qEFzXbtCYAdqiE28UCtoedlgc7RIykySIqpr671EtAQrdC
iebwfTz1H7Sv5dhAGZyrvmI5uOnpVGoFOk2wLnUitJi22NxZBCe2q/yYyAlEeckEXmAzHD30XmES
6HMAT2Ljt4Eil8AUPzn5dg8hdRz6G/q/c3nUQhMZ258wxzyD3z+GP9A341AZjFAjQd2+ImAGdu87
JkawLZ7Cw6LVArl4CafqyWhNvqYXsOgdrfs+wmwys/B/8MLBu0H60r2qSxB6cTzUjSduRGUTxC0e
iueQkQa1A8EaTKXeQe1L86+y8VRY3RldH1Xfos/nK1sAavSKr5VNPMM7ZTOi8+PIGX7V6/xj/zrD
mH9IZ/eezj8wV4MxWX/QfhA4A5lqwl37roeCADqfMIvNwNrt01Kc5J7B1u7sw1CWnOl/TtJpzno8
ZmWOup8zmx85WuLKYvCqOHOO0cUOHNMaMgYyOh1GPzlhKd+Rx0t9pnty5T9MV3GhFBTtxYPIxuL7
g8tFzt2DS6J9E/n3ado0xAGYCuNNUVavd3ySvFYniiHS4E31CrIgiELOYagr5lhQz4sFw37dsEqP
ZeJyIwGdj+xkYf44sd7DK5XqhnxmTABAj+s6nknufNv5yPL/RjM3eMavy8niIVpPksiv4AQs+RGl
HH6OLzV1CIwa8KlmCOSokz5Tc82OUW0vnIeGVRjAv4pFA69WKWDKt0mp4c1tF+/3jxw7myJk9g5k
l+IZK7nIqJ1BCXyPXtMOd5w2ifbM5ndCbATXBExGxnyo9gKFREwCSFdnmtJ9k+CXSwARENDeqjGi
+0bNBHLCh9pgEVeptG7EJua1bsHovQ6F4d6UP376k3x4EJ+Gzpn9vIOaY46Ojaq1J1zxOR/DQGQy
lLebaBCEW8bfMdhuVC7JqeDttD5tYPqA4cor1jX6XymGl6L1rKgoByv76VMWvGAdyZnmZWJWNk8x
0Lfb4TShnmLoR1wS7XqETt0c7KUCemM9EftOD/6rA5Ej6mw+xOT419BCSOraSZXC4+n2prMW5dVh
GRaCWTbeZLPP1znIQP6hMgiDp/Lm5Mo4AC5MjTATyq3bP2jWPFXaKcCXiWHHMkLxfh3GTrfam3bZ
zdP6WsiywMH5pFjQkJnB025ExKMs1a+tonXfwe6Nu1+KEiblr7LvECEOb5yE1O7QaykLomJuYnPw
IO/yt9L1We3zQJGHOlrzbb7hllCARS2xbeC0gammWPVcy3cfaTYXdZ38ew4DKb7upptC1Ffyd6Bm
jVlti3V335BR6oeipDNLEfekfj63o3POoX4zsfyNlt+zIIe2Lh8mBzUzupWuCKejjXFXTK43ptqt
+eE7Uy9ap8+Kcls2qVp/daJEL+qe7BGzQf8jqmkeyXSbY9IgSa9Eyct+pCFUtE1/BzhJY/RQUgRo
mi9hTCVs59mGbzy1AAWEBx/Lwlb5epZTcH4B8J4V+IGGE9KjlwxXOxiYfNb3laiNjSoW8MTI9tY7
v33PkmG4yBJBVnQSmuCQjSvOORA7lL8EBzu6RxNaUqOzkJdro2BZl0/OMAXzr+ADsm+W8r1ZHjZI
+uqLx8Kbb4na2v/xrX6L6nWibS7JhK3WAYk3HzQ6xl/PXm7C9Euv/4ZO4jnQ2PAuPr3MLDPeHkcO
A3aaj6NV2JDuObWLNCdMHdSi0V2MdQcSaO9GqpGEdi3oF3l15wTUxW4nywY30hsQBKL3Q45Qlx5J
9+jU0mt0c3/euwZibr2HzYCtz5PZuNKCCdA1HGqyfgSp2DUHZYUkdjb7n3fS8zCgX5lz4rFyks2a
Pn2C1w2XErBmxG3WuuhcMLkzX6xxnU47iBwc9MgRGNC/1iOQNc/zmx97qE1WJvny+FYHu2X0gGcn
KloIsauRPLIL9dN8+STcTGHEFrUevLYQ+wi6yV4GcmLFDPMaE+Wu4tOmlESTvvXttfRktLSMDV3+
7PvnudvxbvWKqqETf64wBDT15k212Q+OEF8DncRp0otD8BOURyxNj6r8gQEHQKvlob8oTQRQh/j7
YV3+zKf+3LeY/QA7oCcGWVfMysIgZ88gasbgQm/YzsErZEg0uaJiCVToLWeKpTxyFBA6LhGBsF0j
UdeRk2M0A1uBBFqr1XJu7jkXgDT37cBYXk/EMNMzs3+9/Zdyktd9NmzdYIDTW1uWdtnvhSv4t4bu
a06rABYS+L8jqx/cJvM9XJrymMVhSNMqweWPqQFdP3owr8QnTk8d7Ghjkyc/k7DGi1cWyoU8QkzZ
FVj6kFcwOgYUomVWRYJU1bAVwejaHDtXFEeApBOl9n7sU6ZAcClcGF1K/BtWagljbjQOJtoJ4z4J
32r+HVMqe2PSFD9WUF9sC3xN6tfyeAwRDMIGevFmK/wMe3tIjaPRnZpHKnMNzfGqfjCZN3mc7yYl
nKPuFeZ2HyA/rX8klCauaz/fHLZ82KM0JTgj6XOnW6okIyzNEJHOKpl+RTFO9iBE+ZrulwinTYc1
3Pt8xhlnqjf4AYskWX7S2ctpxbVbjsqOeLRSm2SiFBWM6zTXoM10VFwnasa2MqSlLiFoveIakLM0
Y+i5hiPwKoW3IkQSgNiv8yuBozPBaa36zkHYOX4g0vONw6yck6NeQEh2ARMkHsv6/t1/wyfWzLtP
jzXHaXsnQfPOkveq3w5eeEFKRIEbv3l1NiTPfzvo9NL+dMQt9PUwPLBaegmCMC1l020VASdz/eBP
HUFAm9uyUiF6iRQi+VXG63Xah4rIp9stzB3u3RJaCqmErZaTXtmFL1dLwO9Gb0C09bpD6+N4fm0+
NOH4ObsvgyTYF+5t0m8zM5wflr+mst5TbPUzNw8KnNgLrB1fRXq5UzwBqGcD49W5PFtKyA+5jDV7
xwemg2KPDmjBE23w5aU4yjlwXS4I+Sfvg1fpi1ZFL2OPFY50SYZRfe2IVSQ7r5dcXx3ZaQCDnmfQ
uTeuFx9jN/eHrx5iLv9Qa/Ioz6pRvSIREKGfalyhkIjaRzKfRPQUIBDCsMl4iizIQ+dDvqY5aYqs
WWRu7ioul01+g410JZ+ZpYokXYJPRyMAyDbK0ElQxiq7wtmr9/o9gTzhfkeACsY4vs+xRCZ1LpwJ
bd7TtYJs91qD9i8s37Jy3CCqtQP6hZbiKo+8GhtcLsvwHh1rSJS3+q41tK5FVSHnVS35cQn+gTpo
ZW9NJ91tckm3Xm77WSAULl0GaY2qqgR6UClmtdI7kvkOwoxietA7bkwPtKL6w56V40n94NvdCnnD
3VuQP+uTbeHeNWa+goF5EN4ch1qwYMmEHpOuoC02OWwnA22lqw6sBhZIH+y7eXfVo/yK7J6ZneJ/
5Z2KyXbjuAPe9X6+cSsal0D2aeooJ1KsXygh277XLoEUpJQAVRE5ZU5EYajzCZQodymVEq6fAl5W
7kxbUFhNKG8LJ9SytZ4dw577MPJjHn7kjO1KggatQhUYnn/CZ4FU31N0nVh4Z218y9p4IKk5AmwI
+nIOic7xzNbSJms1GQyB7FmAJA2l2TT2DwTIfQUnxAtVErMcizOGOBP6ypVfxivc+NdECqdKjC/X
Tf22W+l+YrK8B2uF05PhLergqN9kYGjgos1TFNGutrh4gtoOaGTLV+eru0vYz97+kTrnQld3RY+M
uwJcnrZVwV8wbzYj54qJnS6pHr4zH156luDOsY2Spb7pTaZiFGxZ0B7g7cgbb6+6HoEKZpxlG3Md
j8oTUHNRNCwPmnLYVDumzo2QcbeuBTorrruTkMLGcONFnqK9o+keomlmFoFtzn4v2NsB2iV+FRBF
WNlVaEA+f134QCsCYssYrGfHmuogYSM5P31LYPKz7EyTU8EZCDh+xmLQFZdSS/kSDsVtHM+ooRUS
6XpmVrx7hNci5mBwY/OXBoVu9VaSmOnoJewZIpIrQP0+ioFv54c7KEqFVqDRLNkjno/qiPKghIw1
crKAa5i8p0Gs63VBLeqmKRCxHwsQ5jU2VF9PYnxdDfxKhrTfzs8kRbIAduPgaiIGUL/ZQv5VlzGn
0ikmceJkXMDoHn5xm42Ymz+EmQO55uaHH9egA53Pza74uewvnqIVHxOHTSD0yBhlbz09Kjmx3XBI
8N4uQL7TQtAOyjC9ORIMaL3CSQgbuEx6ZJ/h3RdSl0xJyche7bTT8lm8ZMSB++IjWFPhqPOowHta
6R23FWkIE6NFuKxBajOO3tVhRrKRyVUGseCVLQkU3/YHoexix9VwmQJ1uPNXPsDhnbmSz35f6FhA
rS+eN/2Ep39UQqeHLV/Wp1D/0agXxt92hnRQEMWOSu1OaoLR5jGrNyIWRL2S8/+5NOGa++tuvBI9
cTxRhbYKApib+WKs82Ms3fAWOOu07GhAYrhUjQqS6BrEqluWZhVjShYV4gAELbV3K8uOnuvQrqa6
ax+jxw9o48mkJI8v4041wvJ1EKZkzjFpnv7IJz05IIyovAHlYVtHoOdeVOoT06Ud8EYEeP8Yorcp
Cr0qmKjTq1ymFxKmmM8t0zW6Eg9D+7SF9Yz8do5qABVeg/tTEcWXkntKtLTm0U6BFi0bcLZWAFcc
b7r3cLoSlxY2wrsPHyPpO9ohkOcRgs6oFABtu7GsYElhxObd7DYxhwT7j/tdjpLf6/RdeEZfUv2S
DLED1PT5rAgJ7ggS3PSY+XPW+QgE6jGu3CYqiPZNv9BYusiMUgiy+1HKT05x6jGY89tktM2I5a65
kMwF73EFdRQd9HBdS4s4KdrG0N44QnAuV+NykV2ffhBZcyJ+R/f9ozDgEfTpoBDvEJc6kC902Xta
RjKaK2I0xJjHcBEbV60Ee1UqVBCqBti+ZmclQ8OjdA4oR3jNI05iWJw7FX5NJYccCKg7WFI/ZeSH
YocoYl9DHaqrNgGuAdTLWYwgIfgOOUr5Qboyr8jO1VIHkQkAGAYAFih878i2Amu090jueivsTYK1
8dGvd4x6Ydq8mHhoTUR8EHBmyMqgmuox5JLFEDh+TMlsB/uNBX5MFnfN5fGF6z7btmnY0VtsNf9u
f+JkmH6ikwRLuKGwX9N8PpBAe9TdrneMJuLMlhTMFNfiAAor5cBQGHvMkjqb8yhm5K6iV5JrY3Da
nJ+nyhP/wpy/YBHG45vL/NU9uy2U7hZkjcYJwrzxGjeSGYvDTkBnLpeIwKjjeW/V0tYexFbG8KKg
c/SQUaDvq7smDYNzHciS2pAA5txLLUk5GfSMZsiRae9jG0A60orEK4SUlIDyGcNlUEkpRdEUXvbl
hYHFjnBct1U4tDCXGEVQUfaXlbY4qzathZFCdPVfPMoAT55dQ9iEoDXADVmYX6SoRthTN4jwAncv
6C8dl0yR+F3OP1oiIHzj5+ULgn3731GLmoJ7NC6WpqAYIu/s8+P/UKPM7wJR/QcUicjLNl7k3a/K
ds882T3P/cf6K61g1QmQXBoTtF9doWFFF1zwLmhcfv9IBPYK4BNrLWu/nJddiY8Uz8E6Suw5CsKI
Men6N2y1+CHU6kukUUDhJ552wtOKpS7VWmt/Xyp7YPN+E0Ke5kWRtslkza9/1DAo9HlpNOMZpMR1
+dh2LUp5CN4I33KkjgSkrHefjeZQ75A5GEs81E99V4Z7yfQ9IhPIp/q/ShqNjBPs2jadep2DaC36
4H85nZPKYl3Wa92lwEetRBzAuJdHfgFDfOOAObf6bil/1WhadTnHW8+n5D1fVlB9SS4gNcTUYCou
F3JFP7X1ooiTQWak8Yu5q6KUAUSod1JrysklWjmq9iP+Z6cYTAhdxKXAaiKXd8ZvX/XbvIIPVwFD
iwIVhzkSHl8Z1V1LZ5AwxiofXgrN9KQeAnDJsx+G0hzWOGAwe//bkoJZwPLns41Mo/azsfzf5zyx
ELtgEXsB4wB4pwmwSZcZx88xrlzBWsp0D5UjLcRBVVcDdw2QRzQjNxxFeNKD8gCmjMUtSEmMaIBp
DUZvTzh5W79P3K31E86/fptdWb2esVUEzNtWSOvGUbb21BhZ+A4dWKCe4gRvkA9h27j7OVu6uXyR
teU69A+wi+O1E1N1EllearY9AX4nbSniKONG1W2ZD2JWrXdfmDi94CkaJfADj4wNoTCP6QWrY4+r
cRzMi6rMGTrw2IyG+Ihu4lSec62MaMNe4zECfWvjXnr9ncCRyjiLx4B4TO7917gL0xUpejsOQMkt
94MXQc6NqqL+788xyU5EC+xHded9KfO+Ula79+ftMitm3SfBOF+kD/zF6G3lSx7dYmhXM5IOZDlO
Sm4dRySNSeGjjNYWqj8PiOSFASp1PO+65oTD7MvBcxONgKOlArCUIZIW1KxPLJLkl57tRlAo3Rrh
nmto1tK9xaa81TRRHw69C56rV4/uB7f8u3O3aY819hRrwaG6TrFDXDLh0icAAIc2QaFvwyd5FZf5
9WL+Y7sXdry6ten2ltDxNZ5KD7zGbVki0TvoG2DvAAbvGBe9zRFv1oM7t5vZsI2Kw0lRUHif3ZXw
YjD79cRB8moYHOw+U4H8jVt4va8RL7bm/56Ial6G9x5cdzhTuPoAT0X6rI2pmfmOfd82szBoEw+G
I+sIjOW+1+9jNz0Cq6b/2ByvJTxJKeFej6bkoY3oZ1zvfmju51eg2wnQgFZQ5+amNwOUr+MxXBa6
hguARjlpM+3Aq90pUtqckKLSKYOU0uxIN1dASxSJWm03jpo8Pc5RDndY5RWVrQRuxUraZ1TgoE8k
TXhkSOcXCCj9vQuMc8Jo4TdqLoS6eXT3uU2B4jLvVD+ZuqG0pGMkDahMdISA+2d/UeP/uYzFnHUd
P6i4W8t1IdgIb+iUmczloihUWh0qGMWzccrQizuVeNFKeAXI5uqq1mFGPb5++jeVbQHaP1V1DZ7W
ZPp6//PJhF0spFPfecRPzxe8XuxTsgPy0kpYTrXIge7R0Cqtx5nXd2jJgBHzpKIPNVHj0caCh9CQ
XiqT9eIBZou61v57/m1Vk0Bnyd1PUuDa7FQYN+qKt4o4qyA16veyI2Kb180zHD5yeApp8q/DY4OQ
ZngCe0cDOL2EB62r7LcHdnmD8sEpKJsZIBEfj//J727MloBsfVHwh1/m4CsPPpH5mChztL4NTCto
NU6ZYAT6nMpdW2xBwFRG61wdRbZ0nty14YTrCjfYytz/7jcomHTobl/CBobh8Bv6x1ot7zCSyx0X
m3D5sAe+cB3zKtOvMCJfsZQIuqUO87Hyf1J4SCzcfRsP9tIk+AEweq0Fqbo90KmmUzyCoB7qUTQh
reGJLA5Q+1RedwnAbA3RZ2e0JFPos9sNB62yTUAXNPiFehkkSnk8l+8m7ShGpeFJtG8QcyqujnTK
VnspaiWvCMr9tNj81hdktiIBmpT0H+9hdLIg42hSkFUTHYQzjHE0CRprMiVV1tr7f6B9Mq1IGhFm
SkOiYPb91WUB2/+Or3w/NAOEohJK2QOf8rbtlG3n6GT+ITDYwtN8fQM+eanJTwB4+M14FtuR/vFL
Y26azpD+WHD78rIOc0nBoQckKf4aMfmwuWKcIsv4JxFmYsUF9/yB6AQ6CekU0aFXyiKIb4NM21KP
1r0zTYWtgMKEUt7n1QTjZy73c+fnjdpjShUwQaWDNydlnrTh35T22PNkYuA4BYjS2EynIJegttgz
sySqIIXSTYR8vTCp8Zcx7e4o1wQ6UR69YYPEols/gZ6pu4nq+pkGgp2oZu4fhB8TlR4uYdkuwd6E
pTw/7B6rQqtb564FQWRW/xnO4+QkXDzKBUHseuxFjfFIJKSU0IZlgkHpcgFIWclAx1+ONt3eiBKI
Dgl91Z6fBz7H9lwoKIejMV/n9B3t/brfbr8Vp7HG30g0REayhDvVucOXrP87w9dvxc7lNIqWdNx1
yAiSfWB+IkJxuk9jOEuEdxu0Z4wK0sB4B4jirZjm6LWrn/h4OA4v+3fpPdTrNdue8sxL4nUAjB21
XH7F6Mpt8uflcfc38h5WE4Yg1kye2y4nGinVr6+lLhno09sob01Gg5bq8QpkRcHDRW33TiKZYbzq
wDXNHeQUL3F4OXvP2zMPqfjf8BIMygeDuDY/1+7AklcT3XWgDJgBeIkGl9DwElm7GZZLu3uPKz0+
muknvz0z7ySspatTRhRLwc+e9WhDfLZekbC+/0A2jFPeA09T7SiuvRtebW0G/x3Qnx8Ve4ONcR4y
nn09HsTPD3swq8JUu0HMid9H+XYC1mBq0jcB6OQO9vomuYVYCmhFXXZRoG7Q7ERh8ZmLgXH75UtR
D23cU4A8mk8/13+vyzuMmLdJXIvgXi/EB46aSrEU5jBldk91fZXvpsB/DSpyha+tOJQLi1qHBtTP
2QFxiksQXWPgY5n1N5mAPq19ozHAeM7Xz7DtoU2PLS1cKKC62Lg8on8+A2F6PzhdDT5IAigVDctl
oxnCPBDTUU/jbl4lAAMzA9VFHagq4lRRAU/fDgOepv1Vyl1zDPXVgzRfA+Kt3qz6i6TuHigSp2X+
K8ifI6vE1PFkOoGMD4OL1PsfxwE3zdj31o6PDS9ZnN1z+mFeKUO1hlXcBKvVTwwRPTPm71//V3En
IAm6L5G2xi0NZHyzz0kBvOTpeGUAuUo8APPRY0X3N9kuqeahFcxGdwGUc+WVgcF3dPcpvsxJS06N
9in1An9c0m28LXo/FUNMsMF9aBzzI9o6ZVA3GZSinKxgH3fBMlZjyaZBCVapGvQlcxDIBRMD5qYM
KewpVgFHYbbUfIRjxuggRYwYlQDUPW4Te0kfIRIryK53aXNqzKEJAxzjbWuO/GxKPxFxT74yRAbY
LLjjvt1JiMvnRrYeCXKo5IdRYxlvOL1KGqYS6m1H7lo4jusp3g4bEv/Llq2dmId+ZGVkzV/37Igu
lEPxLRyEEJeCcGISut8erAVQlkO5XnnmzMZ2PyWSBiciDZOkeBApe6s2mmgmhsRwFIJ3BTc/l9/D
qR5FfAG5AfsG+pixPVvT2QTqyP5tswKryxdE2+xBUgtxHnfpaq53yr52cJs9nhhnS7NkYSRjsULd
JyocsQZYpw55Le/y94GIi6W6kppniBNjlYGXFoXI7JThyvEuT7V1ejyvbbKJ7DDoRbe2xdiymS9x
u+zrCgb4MvRp5EosOqLcIBXscJo+jjyjcqiIpscdTIerad/f0eliVTP82va8aPT6qr4WZjYs8nHo
ksOjFHDT39BOgqPGfk9mn7LVtKiss9bB6cPBgvIXcVW28pOUkrt1P71GchvTAAPTezpaim/tVJ+R
RXzIe6dY+A+xgvBPV1e+O3iM8fJ8TaiExyY7m4gLX0wdoQZtufrmxFMHP+1wp6MeXKIimCxlSX20
ha109gG9Pxap40GFKfgLngo/wwRK2XXgmM0G3yDQ6emDU4px+QtHe4scAEHkOqZUFgSCF79iIJef
yI9BFsukn68cE/Ib7Wynazqej/wUbI+815h8b+RVkJrrCJvjfQpYcN/sRlPBnjUlDO3esfW/k9lC
GQJp5dwbxo9ZIuFoc+sg9HybpDqIOfaulcVBdjSAtYv4E9zo7NrdSjy10o7CDz7jQPUXRbGl2fAV
xkOqdecZuA7pTc+kXlv+BqBMBjyEFhZWaFGOiD9amfGkpSqk142gv79dVfLAY2O2FVi0WCQJdXpl
afMmy17QKCOPKHKYSRTtc1e4FYBWK3D1gTq3mJXv/SVIP91p+il/EZUJb+qIvfTh8nhISi2I3jQi
slN5rmz8KPKQeZ58rmkGqj6gjMifj6kxZnmqHo2bruVV3DN0LWeIKj4RaZlZmJW60ReJAMCGxX1u
j5A4Q+HvEciapMx3bHwKmNGCtvzwVifcEskqE+cpy/G3GZfipmPi8ymldGydcnlDpJASPlo73MZb
M8Io1145cnR11l/J+SeLJp8lMZLzecCtRnXWn2DOjz8HP7WnTz1M+CABjagsb39yQQV4axfbKESq
B8+Ob0zQyfSRnxcxpw2OukRmFabWciYiTjwMymJjpMsSEFCmE4ZS+xfe5rkpginQo2S11yFKuxCV
ofi8hRhzzOraoTx3AHSovYlv+HWxPmJ7xFuBwYgL3oKvpUnwLCVmN5VBPVdVxVCtdck7Fm8+zZu+
DeaDc8iLzXdRyv+xZ2pZBHpJ3Enp3YNwc/OJXp4VH1Yrvkb6BCLuEbx4OtbWpPSQrkUREZiqyZ4u
nAPak6LKs5ndkiPjbZvzLz31LGbaCgY+DPrvZw+V/dxXBzyQpwWr7H6HSmWi73UKydGWlksT4VZw
mQva7Vhcgr4TXTmyAhdkWmze6Am01AOK/fuA25r0m1nmCnSSmUxl+OETUb+30G8jbfo2fkrkF/g9
/SLhTL47ZVhwAxGKwxGIj1L53Knx/iSXkO0JlFUi9XTEezeMXMAI6ooSyuhYBf7MfHSUHmA+876U
AAb5+mKE8eoSWN7Co+G9rWqTRHvF9rcJqnPVsV23GhlYHvFpuglW66iGYmFl+7y0SsSSwsQxQC+C
JQVjD1lD34RQGid1sClmQzPht4TSwzNJ3p8RNqVXKhN0AfoeL/gYHI53KXsj96sPhubSFemMsKOw
JPlGF/AybOyWxfy8Ggni2sEWtcrOw/WJ/zUGBAIFCXKrmgkQeRND0n12d6fTqVsGFxsnDlknDkuO
XBUUttg8IHQO1DFK7ePUTOqJWda23JeGu66T2BImwXduXO3hwWiUq6lov8Ktlg4wikZBtZmTpJQ8
8ETc1uyeo/QD9I/5GCoTSX/u5g9KBumzW0ysJZHdpZ+5UmXC9bai4SncWz3+vv7GGK6D07zet23o
UeLQ4Plj0+nL/cIOnRHxuy5ZiDlVnWYoQoVtW8qx9CnADuBRXa/AzEHRzsgw4g9YLLfZSQ5dOz7I
5oqT8A6UXSN4bb8RQs3qMVZK2Gs0JBQoJr+Qyn86m1x4uA42g9MGX8QTBIwGt20FI0BcID/QJBHq
i72YLJ7kVAU+D9Te/0oZWWDyggk6y/dB7ImbHXu1jTsThlceg31bN81kG+nbMIb7xO60hyKcqy4e
M21rpHXO36yKs2WIJTJA10CrxtMgJqsdJN66tf7CI3bhGWgxqJqswmGLmaPDtcWnscYJ7r4K04t3
/JM5ST3TknoBLKX0q4Zf+3l+3qVzkkl3Vq/TSiHvEAVPA+5Kb+ts4F2kgRcBOslKL0uW9cwXFrlD
biJExAkT66V7/HriY54dUaN3ndZhiApWhOvgvRgNOMwGD82C1nXHxtyAGXtV+m9avb5FGYkvThL0
+M2ZqxhAru4PXZumCaWyTfd3eZiaR+l9ABZFGUBkGqkA2jLSym+HrLhYyfZv+KoGCq0fLGRWlIxU
mcUMH6ZZEYOSkbsRVw8WGOVWCXvQFwYe8+VRsgMa2uIGCCyH5HcGq66Plk8FS1xRxh3B1ugI4SwJ
xMPmfFqnFARojY+cxefYk1prj9Vuh36gpBrqDbzvS+Js+WsTIdt2faddINPZStWB9dA+r3Qgh1CG
hjDygju7/0ioWJTSHaWNJcMc/ksnkyTA7i5XMXGlrJR/5THcqOrZx4ci5hMQAUMAuVateqFo08DI
53Lxx6NKpPUHns+HOB8iExhwyyNwQvYAAHBSd8FVuRRCDk0YAgLGnOqfpyPESsgACr0zAZPsjp5N
QHmD9EPbzD2nUKxV+vSrRz1plLXxtFWFUtMwzlZSJBmXsc/p+BDZvb3VFNQ/z5StzxEfSdHKDvrS
rm+0Yhy7kSLPQOWvlSmwfFqn2aPadtlu9HTRJ5zdJEzN+QOUG6vP3azE/BAz+hBOVvV2mbai/h/b
JSdn27rvb88690EatAKZKtQ/bl9ziKDlJT05FmXwPCDdf7DGgEgCFFX3JWmwUsDRSOTaDXxI2L4A
8Jm9UGF7TXPb/FaIUs42DeSxvQnwbxTQl268/q4z0U/ZXWV8YxeLhzCCpxZe612/f/U88IacaS6G
Z9K7FQPYSO+HGit/U3FHke5zeuYg/uXT5+RNcxDO+EXc0Z7TS+6LdrOxqVGdC0dCVzMHC/n6sIfo
xa+YRnxqteBS/6kywBTaGZeD9ZJnvvCJ/bNq5eb+905MDVtjMXbRuwhMX1d/FQjxC25BMvnuXMxL
U+YlwiXakIBVWV6nlWjRGREaCygH4IXSO7lzxCkfs3K1cbvpQnJ38IK5k+yGRHCFQ+AnUfzneq7T
asf9kLT6NRqYfTt7EelCCGN2LmcKGSluHWV2X47JuaTr7oHrX72waMnedW2KKA+WvGaywOtYPPgA
ajiGB+m+c5W/9gm1sPw9M0pn9OqNtUotvdxzUfhp8paKWhKZoqO0Tp9oRXdZoBVUld4W6JlmiAVG
pbA0q9qG3AOrbTHgNuijvmWdNot9KLoDd3Xvwyw5gz/NUqF/9+puxqqaU3N0r1xI0Jxnhxd6WUt/
HlQu4EeFfkv4MC9ccYmtK6o1gXrdaN6BbWAfOFueoOUTC45+jGVP6z6wxSR7G+ZD9OHZfr2wR3ur
ZdayC0Z5LCy6je57onAG/nlXN64ceED1MOPaWtjyIeFKeqBTFgzHWBXLOjztm8LsAGV+eIwRtxSs
rF+tOIZIUXqIP4duEQX3arLFsMySC4T844eEuSFvW8R8WgMvcRXIcDHs85kVJKV3CSwDElfsJSgs
9VaatP33e7vd7hJc15oyFQs3E8TucKZ3RVD5vta8OuExxamXrjgjP8S34TpP2ba1noeB+j6AtKxt
HjDomRM4A0Cso007SOrOog1WkxEQ2uR9aci2YEQEa5mI2khWgC4PY3pE4tPqnjmC+igh2T7T8C6I
mW3reOe3MiYv7jc+bfHMmmzqTcSzyyfahFkLcJU15UgQGgNQ+hutgesERZKgfXnj7Yw0u8CGsDtl
vqBKA+wlbnnMkTIcPeKSDZY8ARUwUMQcgjaykBq0QzC4iVBHV8habSHclAFZRTJ5rapxORF7A0fH
TTO7aSQa1tP7oIPXFeWj4IKXdFlsxQvADhwOuQFkn8xH1+FSB9CctaSLp5qFKx/RF4EwGx3Qddeo
uaXOI5H5CUg9x8N9p68amWd2egFaau+jNGULJsHUguapMuksOnTXo28ztoHQG8url+jp5QoEhWv4
IOn+0MrgT3vwy4r57IIyzH3wItGSCaeXooBOYWQVqNDFKewz2bw30zvgASl8Q8qnQOYn/VeEmElT
KDubxvJCDVSa5XWiZu0LZ219y6zJ5zmiKvgSGbzqI/dNpjKOrY26hUOUZbL1kIaTrXnrzoKezw8C
srFiY3vHkusl/g+6xaasgmLHD0rVNrcJadJdbyYR3fA4CqWXFyRwpdqDX7oDnlTYwF0JzYPoJegh
Gq1y7UtLeWUhu1i07anxZmodZRarMFfjpPsl0JKWpW5Ixde7aNlgTr1KLLufuCob6aQjhxbsys9u
XPkVCIWvdzH+e3sU2Vz7OnC8XMWbqCx/T3NB881GkPxYbDn8zTqNgVsE3oPerBiwrhq6XtY+s+xQ
3H+0szjjklZqsGnZsLz1oqFBx8oNukX93ZiMtV6p329m9kfFqS64Hk6moR3raBx7YJ0zC97l7F1M
KbIiWkxNZf3g0BOC
`pragma protect end_protected
