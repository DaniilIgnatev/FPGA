
module unsaved (
	clk_clk,
	reset_reset_n,
	clk_0_clk,
	reset_0_reset_n);	

	input		clk_clk;
	input		reset_reset_n;
	input		clk_0_clk;
	input		reset_0_reset_n;
endmodule
