// Copyright (C) 2020 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 20.1std
// ALTERA_TIMESTAMP:Sat Jun  6 14:24:33 PDT 2020
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sM75DpcuGvQcT88J3a+1jCJhZPm2WxOrLHLB68IutjOkOOzLMQk/ddQjxRvR2QRW
n42RnYVCMegZ5NWI8CQVv3D+5M5FKjHiOXQpYfdAZipWSur5oN0rD2j8gplKDStE
lwoiNUOquRAngKHU/wfyFfnxMMtTi36VWcyier3jJ6s=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3104)
p8h0crvsnCGb1C4HA+wjfQksz0Z1rd6CnoyDQHLbLl3tzksDqdqj0KivX9inpZg4
LftG7jlAIqy441khTA2CFU3ck7doVhxiUl5Nsc7kf1/H6aXbayRS3zhZ3bNJdVvZ
9cBnOf/BI/5Yab01Wua2Q2Xss/550kTIO0T4QUGNIeJ84sS8ArOPFAWnezR0OjtD
7AwcnmxsXy/8MdTyusSfRwUrWse3dw4SPO/5n7f1fjCrRoEQdjo8nSMZjji4ZBtd
qCAEv/8CnHuYhUKJy+K53ipDUMFvm+Kd/GhsLq4eOTORSwbWDwnSNE+zeR0T+0ae
ZcXgfd4CgzmRwy/BPV97THpk+bCTKClM09MR3rNyiR7FwbGHk/1UBn+qGH2WdNoj
OwjB77O3pjqeaipTf7rk3B4tsToKH18U4Izqtwdl9XPKm/pKyUcIsZD7DtgrSZOO
6Y3eMGzaWNp2ZgBhFEe9EKDVXhIsZm876IrtQrCxtYoLr+NAr9A5UU+5jeAJgA4t
ErelMDRfOgySauuf6or2/DAot2K9hsBoVAuV/uWVuhnHE13qi5CjrPWdrJE58JOE
A9nTJoK/UWvb0emtkkcvYsWj0yzqWF+oJTqDvcCiWXIFBAzkY4Q7/FJwq7/tue18
+rQhlhWK1097NDjRapIvw70hm7305YcpVErFSPnGJRdg7Zxp0sseojtM8l6urkay
HZvIpz6vOX1d9nFuiQjH0/VE1DZt3E5/XvDGwyoDCpHy5J7KMVlpa+o3QuA9nmk8
VzsBDuxgbk1NhID35U96DrXYmLfttfZVBktzuXmiJEC/Yo1u0bbODvcELggE/N7K
288VokV3+zyXTUbbNDIyEHIPdQlZN6S2vj0u2giT1BnqpMuOGPNpVpweOKnOkhzK
Vhw8rAeaLwJt55HpcbgtBeZWpTA3WEmv15EDb/0HjWmSiaTqnCvzXg/6TX3iI6ZF
ZMx93lTWtJTtxOzm6/8gr5Z8mYhQ/QaipLnsvUg3/qAJxDyL9d7n5swT48qNEr7N
BrtHyxn5xOAaqyPzlrpFNnGVZSjf7DIinSjgWk4jMOmJQSpYNEjr+kqPY8enJ7Aw
LbvbA4Reh0vDuog7+t1zsgUdOvqPqL2BWtAzBPkTSr2/CL8V3aP4Zxbzlfn52k1x
icejEzfDxWDhqp4cOLBO2SsIc8hBy561/ljPYaD1SvcJg8McX//3xt8BbA+M4OOe
i4zklsHFHyk1TXuVMgMwiJNmxXLBH+/LaPvnczggj/Nyll72b8o1CAUsQrow0KyA
Unrc/qozchg6G+FGZT4+2cYt3Nts7r+s7j6SNN/6gsytSEMLKCWk6cXb3hs10gRn
m67Dyx2btJLJ2DVmitUbV+depcpra/Z19XtZf4TRrOUNR+Ttb20VAIOU42lU8LnG
ZQ9F1cwrYdXPnvmjfSIRu7fPYusOBBW60sc8r6NfJANIas4E7mOU4WFhjvQRohHz
ibQDMaBbt+xS4zLup78/VMx2PXVNkRfayhYThiScg6ZqMR0cRF1460OMMq4NWrKR
Z1/JcYLfmou7gG3iOe6GXnoYWViGQNMwnkjJ1P9qhiYj2QXemFUYd6pzX2Yh+eZV
va5euunKh7x3eOkZDmQRzJ52S50290YMJLUmfEPJ7518dg0KJgluf1V2hiHDQ7lJ
56xKfh2feA78R3sRtpq0R+hXKXXxM4ZS2AP+pZOftplonXEmC1730OIYBO6qpSrp
XP0yGIC3+BKVuFIoZ0id7miLiOrCsJa6bmLBB4ZrvRqMH8StGbvSpx8Fo5C+6jK2
b6qfHzp30arKwD6u233tW31LG9C/XCnhKtFaaBWuqHvbq/6P3aeMCPQ1sgVLa8vO
+5EJyDIMShBpx6JlnoPRfuQvZDPvvIrEgswOFYBnA4C8wrIj7Za0C9cZBLHMGi0v
Pjnz0jpgAIrQN8ILsYhck1lsmSAAX8axii4zne67HeWDMd38/jwcd8i2Ke8aT1lC
PJjfbwZqhWl08DW7Klf5N5KtvWf/04mEHI66PGDAy0l+Rlj3OgdU52saeGFuTZ+v
z777qNIIXzCdFWHUdR1sk4DEdfEor7NVABADFk8P6Ebt5/36sOBZJZyvIdTf3hID
vbMlUhBuhHDbEFM9RypiEGzHrKbWe8a867cZPTBtTODdhUb2beILPwbaCxUYVbvn
x6s3x+HGCOxIDgZ0QEly/RVXkLfsBM6XGVhdogPeyvrRIGWjYeqZ21wRo+GXQtwg
9yzON2iv9UTwQICJMJiBlmlJkWMGSxo9aZOvJndtbwD4RRE/N6JPp7jmKB3pLd/y
7XWeP3a44Pnk/E0ijR18pnBiN9V7ibQBdnWSEGI9qrv5CYsN54CMzcVU/X2TQ0WU
beXF9gz+ux+pJryrT4Jx8SgQkaHRCYmuVD27VAqbyqneHYOJxRnjx9J29AUhzO8U
0/HINjTburDN+8n6+alubhp2Y02a8lruQWFSdTwXoS528r3ptavYrhVS9g7h7SLP
M2PfZqRQDNPbTPnRa5gNh9hwnzvzeE9g71d4tacynxSUb//4kSDbbEUMoVV5QDVj
UyCqtSuuPrR0wv4kvprR+cVE1YzV5+DThUp34gnEzYfaLW7aO0ayjuo+fauUkHm6
cCRd44xiCcclW88PILOm3nhGATJME+9Vq9TT6dMcqMBO5c0xhX1tIWOReouYpjXK
rhfQlvPWXJWXCaiBTuGhdD411v05NCrSfflEQAqNl00L5t0uxqZtJqBMts2k2yuK
MXsyaieCZmDF+VRRqybycbU9J9PnqFjQwKvPpeQpbTofOYES8MaYcYfPr1urj706
QQtgcvPa4B4RjIiA6eQ82nslszSd5zcR5w/KhEfT6hj9piPqeqCDhEc2Ng8InnIs
SCnZ36WZfQDzbdSdjp9TDF1mpzusCMzKC123r0nbWoi7WgGPSJa2dOpr4LUQh30B
YqcE26WeFbmLBg/z8cmTRKMjdwWiFJLeZhOyBRZEjiVQW31cBOROMI96ldUYz0/0
ZN7UOfydewsHled6XG+XMaC4F8DVhH1DRLKjECFOJyhLKFx9LKcHZ29Rdh/Pha7Z
dN5P+FkhlWpGEaSZv+XKJKYJ+GcUROJU+ubL9Cs2XHeg7Bvt6IybAwqbS6oIaUsp
v6KyOqqr3bhiYzh/k0zYm2bBKNwQZC5VEQISXoFPqooHw+eKkB+UZrX3HKrKZRww
8eKq/pCfeLsrkRVEOZsED6/A0xKOZi5lZgQn9tt8q2Iie+VPXumvNhvTJ148rhwz
Uhxc79qSV/5sGsYC68540Z9elFOWFU9y4hIQcT/z/0FZOYN5wXd4rKAVTb1GuZZh
Jj28UOzw+bCPcV4bBxUP4g6QpFmZwDwd9A0cJWsBpvD9bN7x/1ULX1t4N89Hn1UQ
ej2y5TJZxiz2EUqQOa0EMXJexas8Fm0RHraSc/FSdvyCOzLDRj2b96ERYl7Qk/nY
/5TeysAudewywZz8FgGoeH8N+F0dq5f/wOU6Ty802a9iL9nEGHVxxVjRzlyaK0Tm
lKi2IBR1dc6ojvH4mha7mQDPHxu6efLSTsmYDqjV14iO3RbiXUL7O969c2MHESp+
rkTjKnqTeN7JcmPimA06h6dmJeiHstBx4sB5McEXzy80LrfQCXRTWNLGuoCU4PYJ
Lx2qGhPDXNva4TZ7EvOWRi1W5Gt7WA2wm95vT5hudy1D2pGHCeC8gg3MxylLvzmj
4hSFFvXbR8hX8fDRC8dOOtGMBETblasAvlcXULN8pb/V5tUTgq1gHO8O9bVo9STh
VQYhc6hJkfZ4i2/4WiLjX1SmSnXd7FVAM1l3i5as9++LPjSoNGeaF7pUnNH/gS8W
Ok9gHedVV1EvGP+TCICcgHn9vqbwxY7kKOcnLCjqSy9lIgecshvvcjsd1zOLMXGq
bxPzJiVDIngZ5+vtYGTy1x5mf9QKeUdEXJto5yqxRj2iKC+ua8QWg1EYwHfAG6QV
ZGYkxHpyM9PCTWYnc5GLOIMnaGgvCs+8IIixpxZn0SDOgLlV7DHml7sR2S6FW1xa
sSPjOx/lJgIcuLlfUltqsS3J0SCv/pfgIaTBnGRt6f4O9R5WfM2GXTGPUEonitI4
wSE5/g1oX9m+QMkgknDz8jh3N94B0EKjmQsh2YuOsNo=
`pragma protect end_protected
