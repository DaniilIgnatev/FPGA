module digits();

logic d[2:0];

assign d[2] = 3'd6;
assign d[1] = 'b11;
assign d[0] = 'b0;

endmodule
