-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ic6i/FnARvnFuzfXPemuqYAnt28LhmPkfQxYAd7TXw9hharrH/Oa3CPRACp7bSX0tDMzJrL6HYzl
8BxoniM30AqvXG0nI5vlSoEFp3yemq5ovTs7tq54DGi3I7ls34ypksBbbBuLqi45rPUC7leFsMYY
Ot7J05RWY0Wceobn6IRDh/8tTmpAklWnoNdnd882XcjAKSIegmPMW3LvqiIS3/dsf1rXqWRTZlok
LB+fOu9iRwn1XigIejxJRjy3rMBmAPVFM5mWK8jdf92oJb0ML+ZVttz/KfW55yQUqy5LbrnmhmCh
mSgT+egj7GCkw+deEgQgcMWTnU3ye0JsPThwqw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5264)
`protect data_block
9CASvLCtsgGRksM6zT4SHgtKxtWaRXndHb5UjeLs1R/b8U+BoW6rQdYdV/38xfntoANofK2Qg8Z2
FqC9zoC0EvV20hi8t1gcw4KKpBZPGwfUtlySrnaNpGDIgXhbYIS1kA/gGSEqLwTHhocIAaNkfvQ4
wrhviFHswBCMkfjROqYmsyHeyVnpGH2CoVMWi3BvKfCxkrZUXhpCOK0hB9zwV6HqgmrB/LizI5Op
7/yoqXMtSKkzHOYp1E3q9Hz+PcQbBnuqgYunizrsywZUkGhXytLWwpcXy/y8hmX+7ke//qNbsrbj
rEAuGfouwWtCOwaE1shNpyQk19Cj9dj46VpbSthUKq72JuDft/tOcfFU1tkIyu38ufFzC7dRwD0z
l+3fFHyX+afLIstqPheYV742fdgnPWZK0xIRp1n6BpuajsYfmFj4HbYXlzSAAQ1bJuCpUY3KiP2B
Vn0nc66FVbcvur3M5rVt5Ctwlz715Aw5A6rBZ8svNTELaisdC5NNKE7e0KVNOY2ySFvk1E/r4+pw
yAhWcgrMMU1HT0NPxYd8RzOH1YND6h7GvTeHYHXh3e3OyYsH8KfL1K9HSq14MkkkXkeqpgcpywl5
pzzIxuywD1UwD6goy+O9vIrCxY12vfgeRmaJahEjJ6yhbu2YBFriWwyfcGoX7fBFsCWCpsqCq871
EdumqtKLpBYX+CAFCUsoCq26qRt03cM36J7xkrVT/+UBMFDIXRm6OACGROV1LLtyR82Sppt+381r
1A99KOpbRVSaQrISl9mNLLTZlLJtCyrppXJDDPrSDyiqoQVyGUQS3Ay2SgVHdtsYbfdEFIBbpdAr
CVeOqcqpXbokVE3QAMk2Vdz7Rtp7sVEs4TqJgbzPrkENhrsUcYSRBO1dmPft9+4RRKyFpkjlwnOT
SAm/Kl/5fQwLSIf+drHq0K/eWdKmvHvVkiOYjiBjzIlN8bYXjJhFEvSjjWVHrhDITFo0emwSs62H
aAYOzu0e78hv6xdMWBb81MFGF+65JOD6f5OTGExy1CzvF9cRefYD3TDgcdEelzqKq8rwAMwmjOHU
aYRjv/5yA4sjz9ysuanfNaOS21ZOy/aNHfslepmM43pzg9RTaH1MovWAruLOGOAfUql+CIosxvMN
rQkTZqjBUeMprQ4hMLM6b0gpOZ6DSrUE48cMckOhF+xAxfEJFdCnPfAxKQfr2Cqwju9SVKUNnQWM
GIuS/EyjZe6MAKdcQrSvipOs1vjB2rOwRRNc9DqukuXHv1/+UnJFRWjzVrmpHwKvqWyXBLcm7GYo
o8SujsaSYJxNxef5urxsIEdsm1l1mBTfsRa1m38x7PrbdMIpyFhqBksOF6XwGOPkUdrRdiOEeExb
fpSzaA4TcqLIkiJw7yqdUjhg5CC9SHqO8Dp8aJF73wn+MuFq9+ir2kE38e5LUw8xUMdMgDkbLkCJ
KJsg6+ZRykSrO3kDMAjAu+1tmb5cAcKul+pdSpfWejYX+9C8hFc7FVEffaliPnY3n/Mgby0YGlBZ
D0mmDOgwd7iDXoXpK+/3gegX0CQxYlSf5RWlGK60SSYEnFzlyTnYXDDt4+RdXv4PIQpDy7HG8E2T
KrhFD0cHpZlDyyRSccXx621f2YDKYQPKOrsAco0YL2gYKwz0OYzUZR3pETwJTFZXbI61x51ZarnX
9UpILymaNVKA17YcpHHf0R+jES2EdSFTIiUWmnzJjGoYUsuRdwRVkTQXVnf9dRLrXqNhOloU/oT/
HZgCXHN4SrhPjPMbMG3uHGxhECFhz68mq5N8pmq+EhGn31Tgp9FZcZ103siK3K+OjPDa/a5R7wnB
MKSQ4M63i+2r3lwptrnqatqE03fyTNenYS9fO404KuWEJ/VcxbI6Xj7h1pzpQB90D6EeamZ3h7C/
Kt/r0qTED53PwB5bFXOrt9r5XkV4Hegq4rwDIkrE8Pj3h8iQ7zL7UR2KrMskbqfJtXRc/Ng41ezL
kCq5Q63frCAOHxOkRqFMIm44INx1OK8gM6XWPKfuWMX4+niXTPHQffGlofHNONeMBSc2V2vTKFYx
u/IfjE+veJYhURiM3//Hivq2snA6AVX3gUbuiXxgx3MMTWtmtxmp+OQKgJxIzAwkzLHuPKWFasv4
5/iIwWjjzWt3gG1dKZc5EuCCA7+XE0mBH6uUMa4zXUKgSYHF/0kgNMP7yUWvSuZcG6RUoEgGSQLv
1Tx5LJ9geVNkuni52g3n8VNcJpveBm5Qt8eGzItR4LJkr454IHyVltyy32YDdxAfOPnJMxwXX7iz
oneHcYiLwtFTs0vok+o+lUG/vOJJ44uvlxKS4DUhUYDwJI/4uL2ZR6JXdVqGY1PrmG6R+xRkvdZ1
qBGVjT+8WbESwUIufqQ0t9AkFT8yOjZExlGqreAim/ef0Iftrav7E7mppglFwDwPo8Oy+OY5UBFb
TnC7rNAQeY/QFnUXImCd6u17jlZ7xkVWb7cXNEAiatr+P9pfU1UuDoM/9KWK2ukE48LNLDVadhFo
YUBgJ+0Pm/BZoaZ0efAQxbTCO//J0efqpdLjpu7Dd+1VEn6Z/oyC1hers1y3PZn7DI9FB4tQW0dI
WyECrt9VJfzPWNXgXieVrMS4PnV+YF/uJyiZZQCRhwOQOY/iZi7mlycq/CKonDskuUO2Gxw01bzY
TTEErAyxdDuUHqtu8828YptkMJ1tNoWClhHy63E7/Cj8sbchZ51pTUl5661hOTJ6lVW9MXNPUX2B
JOD6XcJr+VadNO4aWvPe1wDeCLSCfpG+mH89kjf2oYO9wkkfpTwiyux3BJ1hAt+n9fE3bjMluxOH
MqxlLFmEj2v9USuysbHeUiT7NemGcbgm4na6gXCNgfQDJaUFGrsG1HpW4qLcEkHspXP+29yjO77S
E5gA/cUuaKVm5oF0/EX8zAwcx9FZl9FDT+eYyS0qwuGHOyf08AQMNKvbqLipFPyA3PZUq4cVQuU3
HEYn6hnd6n3U/69l9hngc9nDqE+27sD0kqNNwoxhbjWv1xWbGKrD12t684iYDG82yzclaf3Jb2J9
2Rkm//2uCJ3EhN0HW3aHyG9yx/2u5nNhwGJOiXKBczuMKb8rai40nxQO8rIuTpmloogu5eWLrBFL
MVTbRolQ1iSDM7774sofW87D+rLh8gtQV86tD+/26kKOM0wIjaIk2rAtT5X96oZv5kXsqP5PhJN9
mfsAcXZLtarauzoX0Jb9YFNItUX3+NZRsx6zvPaKIlTXUnoDDvxJaAKz9E1MeL57hmeuZBLVlIgN
fN235YvB7od+m4GhiRT816ux6JCSJa9rQZ22aKAbb0d5oPpaZZm8YW8D3ce58A41L8R8EJ9p6a6Y
Qt0VIendMGvUSrYklWnV5PcjO3kxgtPSxUwQY5nALpmIWxFC9HFcLj/KFqVwXvutQhBudFK1Z7EY
Yb3IJ1tidLZWsQ4MLaa+TweZ3sG8ECEuqbsDZJ7aP+UuucRJsk3olfa0TqTpTG+HayWm6QM8y6q/
CreD1f/PJCnqyaqlcvG8/hXCKEmw2NTk6Z6yb6h2hY0hUxNTWlxN37I2Dn2qfNdx8AulzgIjjT1Y
CrYrvo3qGQHMgt8rrZv/d/VLVBJ/YXV1Y9+456eYmNKZB/PVyV2AlhuWqUbfokFgVqTr89kusGl+
NVjcuAH9F85DuW80Kx3AHqWOJM86g10EkfF/iIg64/T5Tw8ylRanebwAGa7D4/jpbn/mThKo+jtI
6mK9UnyZa1a/AESvhpppAkbbzpotKdCEwxDefnlcsL9FzOKmkkjwCbGSIYIQeaY8HN0DLgTh78C/
aXmIshCDSEmYGNio4weo56IXax7ZCQ9INcxTxvZnpsuYgCyVb2XJ+NUYn0teoWM8TTgI9zF23+RS
kOux/d0OcKwNcDiJpAyw4dokX3NMxINjqaqsogBM686vGYM8Mc3zQfz5ekqlVLLg1iqnewQ9tGfi
gK65tb+A1U3i4+dxq336PnrrR9uVyMqwOUaE0sg1bmEH7VTeE1mzKKyF/zZv1Q1xqB/I/C+WvnxN
LPvJLiMgf2Ergy/o2rOElNbZ/Z8GQa4V2S18oO6PfUjugW3Zrv9+JTb/XFBGM0C5Hm1+ILvakTyW
VAQsKYEmah1MfBLJ5fS4juDVKj5YQ6oqgcGELAhx2mkcotd1S+664zmkNShRGb7fPNLudCnOSMh6
uMcyvKHtZVntfmxRxCpqzR8Ywn7qnTVzjrsjh/ijdCECFt99bqSecyaa011CTJHU09C/SFRFaJWj
hSZkQ4UY4kw1v5jEZa8nbcF6gkGX2ORlgvu7u/VsF7dDGFGakW6fs+wimCIJQNL1UtwN+7Vk/M8N
UEf+vVR59MzaAtNPDJheo7eVHwN+XioImpJS3LviSvrTA/WWuG3aFuOETAuyKBRIEWB2LDWTXHLz
daE3zovnFIbq2ZzOM+iitrINBR9YuLCTavPliWlSlPs6KhIyTneSigHkoNirBs2ZC1wnPi9Bk7WD
v8K/JO2QOjw8LNxZgG7EPWZ2vhDZDyBCqh/csbjpo0hE66WD2pHSJjAp8d7ArqJSUxJluRXGXU9C
0UEjcYdGM6AvU/8Xs10Tk+SQqsU/h/wmOfF0PgKGXYrXbcGEn/eC40CHNRYTAZMHC02VVL2pFpV7
vONIOK6ECvEWhder2flTKeAq7tV4HrJuzXP8md4eMmFB5RYNfnWE8XXx5whKUnkyxv0/2sxzM3J4
7dA58piZ0T+6DPVgNMYRVE4mp7UUSHdgDCbkb7tGiagROstyfanE+i/obC22GvvW0fP8pGtdfcdi
j5BsDgPxWdm99aoZCcf/sQGVsM3ER/DZ15Auhd+0iPCwoiWzWas4QOIDIEiMqJnMY7Rf0h1C05At
8kNRsn36dzoOyehiQnxuOzD4qxk2L2w0gE5t8AmvRK2dT+lZFaV49sBcfia7YWrrGDN/Li34aXs4
3RHR6shfXCNHiMmzk0rrvRTUnQpBNfUvsefdlbC5awhFcf8bA9DirENaKB1Dm4/NHpk3m93kisiq
nd9eF37+150PtfMCisS37lfn9/MMQe4e8rxw/XjShcL2/imFtz5T3sf3bfRCJdk08GgCF6jLX5/D
SPne0h5AotzRwVkaG0t7kjqxH1tQ4hU6d31JwsdEF12YLpjAioG8z/es3ePEP3nLp4dPrx0qJqE8
3ZkpZYp0WTP9zgJ6rNP0l8pVGgHBFH4Hn4vNw0o6E5SMLku/hotGdtRlbvOas6GkTmITCoqNotGq
cTW8buV4jjow3Bm9Lhfq9pNdsaUFJST2Q0k3ZASixIfVAdPFXnbddfEE+s1V8vMOUgwEp2Qs1W/n
k4NtsaVl/c0qMsvxWSL9QU/tbqXgnWAuyQlBxZR9cQ2H0MFRmN/2wboYZWfXpHJONEQ/aQTku/Ci
jfDcd5NoeMCN1OnWXSpKcYGWmZKvScvnOHuR4P48nEOiof5eLV1LDPltEYe69wAkBmGGjOux4jH5
1n5V7vt1jsIkgDpNacPKRwYbgzaXmSbzaWaQERxA8JZMLFC9qPhmAEG7qaB82R/leFASqnzL1U/m
uSSeV3JweoR8FhQB8L4YvoMoqb8eKbf/bphVxPe+nC79NMaPHc6q1WfaxaMGB/krLpX++dvsfhu4
+DlPQ3r7eNEAYMVnwjV+nC3HMr6E/Oh4P7pvaUdEnoZ+O3hHOn8PjrEjCBZ6eun/1+Z2Anc8Y82S
FLlTLgp4FYl6SoEk0IzbdOOPyiYHH1bw15x7Lf0NaN7Ja67XGVehIGaKZiIW/sXQYz/um4wbJRQG
Ydc4ZlIqMiNB2jAYOUZmiivimOnTWCJKKzCDNN5TAC/F7F0NaiHKTJeZTdnPv99y4Vfnp1r/61el
SrGPZQsxt8QPIaBSLY4SHudnf4cSiUE11CvArJ3XBllDPMv1gs/nrcvV6MxtBjFHtFUs2AZg4c+d
i+CBmzdLK5/rJpP90HqIARzDSB+RLdscwihJenPU8w9bLQdMGlK8H14QQ4GhfSmp6WiNkQ1qtf0A
CBou8qNLJbGWCETCXwYfx2N74Zj2ab07rTx9L1Q166zsjWY/uJNqpHRbvpVz3F9vaofMc+5aPs88
1LyV7Lill7VZ+Gatk4R0K153DL4KY5uwbERtT4GogfFwzitppfvDfWoQYYUJEsndrO6eD9zPW4YX
VHYmNoU8/aLvjYOiWxYpo4bAwZtOF3cab11bEPjXoQTjUdwflAyMMVM8Ifa3gAlB20WwAgkqXpxd
62a54TKG4hVklwChNk3xHspTlvlb/cOX99/DzFjMqbP98nJgMnO/8L6FQ7qO/JkfA15hioimr5/j
SQCkVINiWum/UxsLRX1cVTqSCK5xq3QioFNAxlPvend6oDLrvXk3t46YtgU96nVszWB5UrwXc8sq
tzWTfv/nRb6/apYVUHq0NYMn02PHplEfnIiLWOJWU1gPbEGIOzwfo/nPFhey5sE79Q8nRuD+j/GG
ytGYpjw92qMQ9trj450SA+JE304aZ6XBTgn3U7YmaI3ASvaBhRXVzZ9tiXtZqgZe743fas55IlGo
fY3qnumSR6Wsn1dE8og8n9ybllbSWn6J9R4EiUY/X5ntWfYQgRpzXpQv1kpB2uEUc3kuUPatqa31
tlXsB6NnFEcUjEr6qFWVQ/AKhpXiFwE9ujc1OxbkMZxEtgtWIWtnkUyBM0c5O/7EFTfQiI+LtjDz
DmAoSJJ0KsGq8e6eoWGj7B6cGR337icVIlu0d3n7MeHsntgBwXNlsYG8vfrt2lSdNTI3dvgj/ZrE
kk3sojIvdTzItihHITd7ybTRvyDBv/c2M8IZNmCD8KNi2Evoolu72AUs1lyBF7ttSDt+Z9rG3Ss3
0V/8Sjw52x6MrrsPGw5KV/f2WpuTjyscTmNEHVGv6ufDOk0fk/jqkzwwe8YoCROana9XlZUxQiRx
y6vj2u/0NMrVLBneSLNDGvDo0lb0eO4c5cy77SuLQxHhr7DIX/1S28hHNl7ucl4NsmP9QNSf4nnQ
UsxFMnB/gjSaZVR1u7FI2OIyo+8=
`protect end_protected
