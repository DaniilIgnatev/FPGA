-- (C) 2001-2020 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files from any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel FPGA IP License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 20.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Qc1JIkO81F1th8LWvvNLv1PePq07aoFrfdnE8w3g49nSr55Nt29zQgLDy31x9v1SVYmY08uvuiqA
Qp3uy8q6AoqvBDt1V7lMVJrTGdFoT51MFrYtmdXL+zrupFkzUX9LG21ygYF0JwpUrYcOEayDMkuD
HssYX3Tj0qqutF3sc9X5pfQ//w1qM5kVzPabhoQhE6f404+w9kDmzgL4WmeWF4Y0j9s+jXLKjZfU
NeJgIhE9wzgVkqZ9Jq/ho9/E5vIeof0zl35+iuBHAu+TETnZ7CUKKwL5oqE6N09ckHbgkaJGqP5s
xwxhAS6GWRcToN5PDJ2KvqBp3zeZkd9vwZ4k4A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8048)
`protect data_block
u1ZtKJir1mN0foiG5OgY78WAqeDIqxd8uxRDKGj2S8A5ECydxonPUGLqXmbLX+UD9kQccLYP5auY
qrym+OKu+MqFjh+PHGoykdzXmlylkR76IDoHjuWG7WiRaPuTsj8aSzVsic1zQRVh1o9NdHOoEvc2
UGUrnnodLSaOM9ebGFiwBmzczB9RLpwGCyOphViSQ0RXuSCKpKl+vEVu4l5B0UdiTV0eTYeuixst
IKUWKN/8zs8yPMN3PkWwGwiIAJeqluWyA4cWdnwS3yvw2z1ZOzTjsiPB9o4EN23AA0fg3s/YH0Nn
YcyEohHSCz42R4vMgbCUC8uWD0RvL/5eai0pEkl4tEOblVkma/1LPns50XElrNSyocDnUy0MdgjE
hqggf050F4OqPSd2Sy2uBzFyawbRIx3r9V62pASlw9pHMz47gFLl77XiUCExjwQ4fxssOs2eKzps
qYAqRfQmQIC5UCLL/ba9Jv1rLbl8qEXXFtC8VXQbs5dz4umynU3I2iddxPg3BGF8S60QTltVqGXx
TaWZ1FAutMpLIWrcKHuIkbVY4Y/Mp2EZs0stit5HyCTVmerxMqtyfd56w6YFK6eXXE5PMA5eXdRO
oYrNA5cEIoh7Ha7Ol0zH+LHywaCQxUo5zxuspDogeP5Rok3TAoDNbV2xVEQRfMq/WnxkIKV6TMEz
h3mJlhhrbTtVVMtadCR1B48FeDxKUdiugfNP8vZ1oIQFBQ834Axv8zKsJCQs1lJFsQPA3NPBS7mx
G0UiL7tNfvYz/ApW2M9Jhb8s9QFJge3UEJQNI9qKScHx1bqojnG+/6Mixy6nNN1noZZ+8zTeXYDT
wZedRYqY5DFMuFAnBfDDlXE8iGcR1kkdQZRXwrMK6+BVbPYhyMIUoeqS2IpFuRXl9DerGaDH3H6e
rk3wHFEOX/VdbAyqCCdELMmuiF7XDvL147zJd8NVuWwRWdJTD6Wi2BD/Gc9ZlktKcx2T70OilesO
nPQWOKpVtb+JIdKwVvL+TbA6sNeLL1A2E4eaXbIWJBarTgdaJWPaSXrBPuMDSvNUYH/J98PSJ7/l
FUnVitVo6LoTHUEwVV9nZ1IPwBOjZYT+UJGCrCGmjEMyzTxM2WzjS059EssODPElArBqFF1TvTkb
+MLMH7nmVw6tjocW+2e+WgdLmfLuYDHl6bAj6S4VMDxkXCBajtMuEGQ1bJO9ocjTcBkScmo7tMX+
orNb1vSbDiU5OAlkTVXqWyuyAqQ38eYjMKT9DtTi3rVNAVyi/6VRmp3KD5pyTVzHH5M0P7OkowNM
0/+NY2lxpJHuOQwVmQnVJTT0SxTQekV9MlSj+w6MoJ6T2TeHYdf+mR7bwQBpVwZBsytCl6hsExM5
1tvj9mh3nqhWTpL9+XAlPE1eS4jk8EWUf5f5b6X50pJXk7KDlo4uLuS9i7oGpN1XiedGHltTTdQG
NLhFHMldmPYK6TpZNSRyQ6YneAxkT+Op6sZQHJdL84fYEAxTN6yHbfzLgWVCYXWBjzAm+PO1vyfz
K7fgB9rEoOOTSAHMTgQ+yZ88AQp4GqcHV+5u1dO61goxC5iBe5S2z8SzJP0bbUc5+Q7Hzlds+ydP
tJjHFk+EyGiuC97DeF/dREqd8D01etA7+0/oKNeqpti+qgYytoP+LM9IvRbxmBN1vRFnlbLqomqV
zky9ZQs/Z2NwRCA/mjSvEja1Kejr69+6LPo/g80WihfDH4NxKRR6fex5gwRscmABR+JHZkE6QCe8
9x+fIrEqU5K5NyBDYdazrUnV+8bXDjBigydvesmftOn3+BLrHtEwnSjUDzs73WVpFhWgQQORu8ec
SN0ZLnyWoBeZxyGE39SwRe9xXxrcJgGiCa4R2ZAGok678nZsS23lE5PdKjqJbgtG5+UcyPQj32gy
27lVcaDU9IB5p/VHRksw+JOSnYU+a3HUEcBCE2WqecLtAwlQ+LLWbC91iflFqktxZm6oSJgb+LtT
6KnO86FVHXj7JiWmzz1D7dZDWKqatrj3dMqxgskk851Os7ZRrZE3KAUaQx1S1N+3zoNXjv8FqrbN
Q31I4zVarUFz7HaYqsrc0Xv3nzNm/mY4rGOnUCJBkrSTe52UXSAKIMYkaUN97dFjlYarccMGbs8D
47XKU8ohhdTr35QVrjEP+K3xX4IpycCCmai13XSGtkYVFjfLVs6Q2xhdHjS/RZuNf9gEY0iBl9bU
ugHldAiJKJveZ0VYJp0y+Opvb8CSBTBy/bp15qyWhDcFH1pwxHauVRdiTtejdJ6fQ/e3pjoM9yK6
MQPMYdg++p6PCoUFLhCpbbB/XugUq3FruROknMS94w/5mEl3lpysVJAbW6ZL093KzMKXn1DYkXZo
FndKJOqOKFSc5lAZgoCcQqmr6Rbz3hxOHa+x0/V0/z8mT66A6ZosdOi++plJm1I6kZV25WxxiOXJ
9dD1jKqTMw82BkEnUkdjDSULEKkhdr+KVzy5VOGLo2FhKsIuIAz31XgINk/h3f/xacrTlBleJkdH
R6DfhajF9hF+gl6gDwkXu08REUeRHa6VMH65HXtGUgOMWD19XvLbgA1FrTpaW+ULce5PGzthQY6w
q1JC1p7vI8kwiq2z7R3kIh7k48n3ipG5VlO9LI8QLYmB+xX/uKdXwl4unUHFMn5cr22P2h/kPfeD
YDzaO15bqt7Hi+MAVvrWGhqK91D5YSfwz7iTPsY8C5TJBydzWBrgDISJ6sX2213CamY1zn0n3zbW
XlJWChqzNNKbAi8HaBtVyjBiQcUtdIwUtSc745ony3bXCTpPn/a9NPVToYaUS//6clL1L69SrsiO
bAmyE8j6v5uXI6OEs5I8eNj/MHOBc+YlxlrWqTQ30HBBzz+n9HfcteTTgeuzmACS1RTd/eGxcgJX
PTPtc04UZYvRUF6LZ73C0T3Wpq+Kc97RwsdauxHS4xCBoOL1bvqQvf6i1mBjWAoXqMCiMempMHqt
qL+M43Nj0IJWogeS28Tjb0PoewFHae21ZBq0FZ/rdxbst+ORsx1Pmzj23UJLau1sSuxe1VhQWjk4
F6kYBcax4SRXnDmP4g12zOCpbGX5eHBd78OUK9N0yR75Tta94iR1x3SUznCIxa7ZlWf5/QXYEi5C
K3bfYSzpWsQzer9geeg34zXPHdbTN2jTXDSTXmgsyVF2i5I7XmD/R1ovxu7TJ7RrfPl/X0sRooAW
BOojTw44ONHVj5YuEtg/VqkB5LUE6L/CfqvdURKI2mxFZkUH9jH39cZ+Lvh8tMEgYuidCrVFoCkW
pUOH+ZJnaU368TgsOlNgbyW5OIYfj2OXzylGgdJujAaJUvfsfdSi59hxltjaAgDhR6hIrUfivzHf
HSoQ9/YKv4uF+pVL30TGnXPTerHAgbELJf6aN+V5YkvymgemMvjRm2NZoCYbKS5WmyrUn3x/B0Mu
YdoddkH0KBfTvXnPnDnRYRnJhE2A1Ctp17ZDy48AeuSOBzaQJprsZzJr3b1faq07l25tzkMmJlJq
vcMqyW5HvqIvTeeDZbThGqqR4cyDa6VXedU7JHKyrJo5t55eWA/nR5uvgjUFoW9WGdXn5VcNYX4u
Ro0lEuz7hj03/D1710GXlyXTxQsHTwVT6UM3tK811DFA53PnuHglQQEOA1H3+Ez3l/54cdNdIG03
2Cacd9O5971VMQr+G4suCUAWvAvHrQtarG8adq7H2piEqhssEyYTvYieMIy4a8sd840zSqnq6CRy
NHzIFXKOOb5sQQHoP0VaFBTDHAjZe54zcTgq37L6SY8ALsRWMDf6PAPn3pZnjoYvWo4p8qJkXSJC
qFIGIMlCUjPtrfXCOdd1R2ExANu4xf556aEDQxSUE4I01BJsBitad00Aht6oLxGNmFNzaRZq4fw/
C3soeB4YIsBxcyS9mw3UKd3aavncyFvA3cNgQSRT9ww4PSrvFoiBoLcWO3+i6UsIXxUaM40bmmpG
0kDYQRMrej88G72o4W8+Q1e5ge6zakFCQ2FAX/r9VxW3Zn9uqTI86KzgPoxikBW24Gyj/oF3AYX7
UNukhhxQXknIRobKAgBZEKvoABdUrikUdym0SnJ1i6b3SRNuFpHhQdGT9t7zkn6615mEH7r4VdmJ
1NlzTOcqlyB1/PoaPsa0Mme34yu3nMZnhuIRqrrgmYSu++Nky7lCVnPSfcBj40l8MGWQA+j4V8Zp
WlMElbWCofTJVbktIWz4Cg2Zw6wobyZvY7hhtKAFnge9UfoInT/Nsjckek4duGdfD2rOCjW63KSz
1+E04a9L4Qowmoh60f62zW9zSVq6Ney6hTZeEQcHuRGzc+oVTWthz0g42Yc+ViEndaMmxv24qOem
kP1PFIA1+kjM/fXdt1haILG4U6beEDREBrVSw96xeTCEzUABiHggK8gN6hzdc5c7hrib1gXjyLio
Wk/hd3SrAbkjsFcRlLnQpTOd/3rjtzzEWqh565NRw5m8E4Tp7r7aDketVHd2yvJPkUC/3BjVg4kh
WQP40gbBf5meyTLAdYWdgoKSTRAoxgBqhbWHSxJ/ab6zfaiZCWvmKWYL6/QZS2BW+W3i8YNH1mIi
jhl5ZVhiOF+X+DMuin7woJEQGPgZNYFJk1WrNbA8Nvdq24EcywpIOlm46Yx9rMA7BsWGA+bMHJH4
rjJjRrLOSxNhqKNFAxkkXd5Op7CSGn/eQPYOlLqwHdBhtdiKuWhs9P1ntaB9/lwYM9hlmbBUavom
QvgK+ZLV3TQJTPq3gOpofbuCxfvsUk5Nb3vg6+jX8/ELSjrhX3TCAhOnK+ctc2cY4nDoxgQ6kNaP
ZlhK3TMFWv0lZtuftImHZzIIO5w1U9CstopE+1g4CRrGN1bCCZY6O9FvVcZxgVFw67KgEJJk8xOy
XI1QwSsdo/HExhrmHhm9Eko3FgdTizBRNYfrFeo0g5rmaCXK2a+PKOeOfMbJO8i0lpQTW/OrS4Ef
tqexUahh5Dyu6hScsLsNvFDn0FhOBKiAElvLTaG5jJ49KP5GAea6lxQkr4Gb9EApMTbIV+JfSD9T
Ansmk52OJXsDnjHBEaVuFR0sIQr6sCXlZkJJC75mR14HpFtoHgJ/rUJWH+Z9yrhHzWjovGnC/nJD
wxS6zv7HGclAbScP7w+RR6lPM8BzFSZyD3DN4tV45jbgKhDcFQSJi2jgGgQNZtNiw+MKEldNkmZW
qvaWvmVeDtPwlTJMNxvQap1Il5U49owjv67O6zfWlH0o075555emiWeBOR2ZJ1/BhKTsxgpUtoFl
phqVLMiKPlsSbAX9QQHcFl30RqG5ci8VeQK6cK+rrICwBFOX+m9btqmhp7qorf86Ft5PpDyr04uR
7YxcszNI7hWVt6cO/FeT3fLGcy06a8N0L2vxmfRiPO950cekZ1u5u65Bur5ltt8eJC0Xqn0WXtLp
i+kOeuMcA5Soo0Eb/mRLoU4rO/sY6tqOggfvrQzbVS3kOHg2ww0/ZpYNbfJgDYE+LTN2GHVkBVMr
6U2fgmkjmUG4GPEcKV4SI5rxYjkIGFLadBUm9x4PqhHhiOzjWL0D1SzoarKQ89/8510a89Kjdsxw
q7Y/Ohz9XWAZVjvFOG3O1PAKTicB3lRAdclMUgEMjbyCKmj/RjT9NQLkY9gCiYJLmAF6SGQ0oLVQ
pYKcMHiQYEmhtKOp+FxvqrlHfZ7hnZSLX3ZGmajcJWx/kpgnwwu3PWcwq4LVXmx/pVZ0AeBhSeOz
1nUI4JOVb3vUhd3qz1gKI87gkMfE+QQC1alylTKS3k8N/YsNXr1h5j2j+RisIQXM84SqU+t5/tht
MBvirNI7Mb/q/vdixCWKYeUVLi4bXmftUxuUsQVeB5DgI8lEyMpZQ6rl25U1Ml3S5p8CMU4PYYhA
Suh46FY6MxgOPKsH8csXN2vuoOpDHYp/WwocVxRqhvtBEz6DqMmm1zjzQoWYqc5FBagHrEoPEvyE
SbalBCbByHkk6x/zYz9aRMssttry78pb1PE9/DQOZUqoy3GjRlypT0Q3DL+2jryXeRK+LElrU6Kl
Pf9uN12MyUd3Wgc7EZbBuKqIMQEYeIUVHCO8OdTAOSSiWRDuhk97oia8LvnYeu1D3ObX5gn5KrVe
RvPO6fgKhOo/8av4JftEObFe+72KBbOi9uMz5meYGn6EcJDJRxM4iX1Nj0rvuacUgnCbl1XSf+aD
s6/jYJGuBhvjwvw8sHfJ50KduA2WA/AczYKyzvnbpnEA27IDnMj/F9D0O49CDh75B2Aq6/cDn+AF
Z9LQCvrXUTVA9d35jfjyXsS8jIK2DrCoXNpjrsM+1HAVrb/uU7nlc1Y236c5BjEZ1SkfhTQ1aowd
9XXMV6l0lEHolAYSg7RW8kCS6PQtTKRYHfxN2/97rlTB58kWQdBwkGB/3mLfjtL6xRMw7Ju84I4j
5b8rhipCF8OFywrnRgirrgv1e0ChwyRb2QrPe8dTPidnDlriiS4sSGAEehnQ+0bSn03fQ6wBj+Z5
lryfiGAA2Jt3o62i4zuKZEN1tDRb56qUpUNwzH/sOtf8cup/Su3nOM15OWoyvqIucHIu6+NKb3WF
9NR1Wp4E//Itz9vFzXsydxJb+vViDaZL5M1sjj2BdPBvlsQfgEobZz4+2LlwOHKh5BOm2pEuSaN4
ekm0goG97RLTEbUoy4k6XOAtHDTNERFw84pSCuIlpEVtzv7o3tDqJvV/MYzKicDiHL87nIgT04Ct
/8Bhd6nDr9Wwbr07pWlXuxkxW91RUinIodKwCg0HZVycvqLHX1rZenGcOSiqXztvVrm5DaEFPL83
uExaNxXTnAt3rVUBJz0O2uwrVaNsCv7wtC0Da2hS3biqJOcYwxDEySbcsfQT87pxg+2HEP4ZOXck
lKtzHAk16BuAOtb5G0i0RdpoW8Fdh3VCPyKEJJNPz0YRF/MbT3QC/Hy2EOKbfi5mGcQPIgMPfPGm
ZMMgGdk4hE5v44yy8+bPezRnmZjucosfuKSKim7g3fEKv7aWHsI0fUqcce83h9ec+FZ8p79QRCYC
Sht+jiGBzQqzED+X+cYFbUy66GWN+sv8ImpNAHNxTTYC1kxLzlR+wQPT5dqQMBK51U3+R1Iacwfc
AEViSsMvChO9G1ZNI9hJQukAUZ5+htzGpgWSMpDpkt1VYErWsdzGZnTN1/fV5rKETXfzcsPERQ4Q
kxIJySrXjFpAT9vEK1sTaV4sdq0ZAVa22eKZQDV32M4ynLih+tUlLmfBhR5XW5bFjrA1uIeJQIoH
424ScLVsLY5sK8Y85nGiPoQRD+jXXh8PIbgUdPAGXSojeRNQO7nKUUmcGktvb6aoAOuQ4BsW7ci4
SYjT+O/J1Of9qnadtxa35Djxk8SS4C6dv965opffQA67b8tE+h3gUzJnT+Fnaj1BpAtmyjluPbZ2
aWZEPjwGxVC06VMK8JPBj4W6E9p9DecFdSaglMvab0lvUR31G6hSxYG6pWkLxhLXMIHhcXJIIifP
hq+S9MGjX9qucGC7qBCF3HfUqEHqcPCOnSXjX5GMcX+GppyWOWiPwZRuwjWhL8TsZp1AMa/jcYIo
9chIoTHos04k+vdT1W1aRZaQI9rq+V3DPSaz70C1Mwh5ENrzdLgMO88QTxwxzcwQyL5HUegR/tOR
o2RcGaiK8ADZjD1jyJolggwruNLD2aLI5RKHTqJLy7IkOnxdMUT7cKLgTQBjkdkUiLSGh5jp06Cq
6XIxJL0axDh1xVcVFkzQ5+TeOlKTqh4CpmqtGLrf/9O6VX1ax18wo7veVnaqSLftvfHBZ1VwkFEZ
JkuIesM4iZZg+F3A8NwA4jQTYO21NrsBYb0yHtJE3HVhLLoRYcQaOcVJgOvSD8qqEvssi+dF2Evn
UzRcXwok8b59OQrWo3/olwqFmL5CkQ8InD60nPnw4562ubK+Hzwzk3Amyp13je62BNMcz16XSLN2
0c+kfCW65PPZ8gW58jbAACh8wYm3qWMudWF/aMQ9q+7f1aShF5UwoSFGd9xZbNXiRTP2uzgzEIQd
PNv/MBqeKHrL+Q89qobaQ6alyaSTk0hdt28Qnej+fQRC6wqQ6WzAFkIwxFteTCKoq4d6zw35M4UO
AY5hvv7rhJGKdwGcWGU2G4MIWh0Kv4qHF1J1vX60zmWctY/DbD6BRHFHv0BusS8cHjRtg0OIZQC7
xlqWwC8xD5hHSG8vtYnAQ/Isv6gFJTQRQXDltkipbKkN5L3PWY88hOlYDx4X5Jg6UATYKxCXznBa
ZQXtSuF5ljheoc7ktwhrxy/6dNhX46DjYAEqMWgWkljNbXwrOkKdHD0jObT1MxmY4VJE8evBX9zC
EdoVljJISa8g6tpUybanxLAKoci1OJRGEMp82YDNFz0ZtVzT7LwVdoDpd1qjSKGyiLIZQTNWeouN
qYYZJjqLQX+cFLfALqS32bJYFtJJ4TQPLsigk8AbrY2IfDdLaxwYsMeaDyM9ptAkrbnjhoVtuNkb
iNhmt3P0CiBBewstIHwV3wpRkXBUX66Jc9FwNvvsoDOMJtXBG6/0Jzcebk0T0ihV6plkvjjj9olP
ZIIdLpKrt72KQ9Ob+KD+J7Qg/MVb27/dUMwu4p8ohg+Cl6tv3GDFrMo4EFK38D05mZDQxhEfw2ns
THJ6CJXymd8FUEhEIQnh14Rf60/L37qbsFBbHNtrXwj6+fyF2qDyDAi24uI3TobovDTxirWHUdwI
w9Tq7B0+srEHsiVH8OMY3/CevOYJPrZZZgHrC78NoIw+sm5oV8FfAt1psQeLJN37TKZUKV4IPUpC
XfwuZ9dfx6zpjD/E6l/+3zwCz7tUUj+lgCLT+W45n8B5eS/ODeDfa0lQY3Q1usmjVUWxNZPmoW3/
+4GwNHw5jL6HA5wvJPhVUuli+FfE/yXvUhUoM9j73vpd5Z1ReSVpp2gzvkW0zzwwPfs2bGqATQvR
TkkXEB0XhP6eAH7ir/22+bQAcPXtd5vqCEbBhmP6o+Y+uILIyM8sCKZC9QQT75tD8xzPowJZyklZ
g18pULe8c9jMTtMzsSOZ68Fi2oYha8KPi0QzTzHjWTOWbXjAYsOUsobG/NzoSKYYfMGOK048iCmI
x7VD3e7Hv5L/ujopXQ+cSw7Ujpy4II/o0exEi8xstPnZVEYB1o2SU4MrW2caTcqL/IrqVjq3Twg8
YXXlVBDLOyMbbv6zNi2XPKTEmSuAE7lSvmgBuWXjvhTYTGOzGesFEqCRiw03NkTFhGso0LqKSCW1
pBkBsIoRE+prybeMAQOtCvIY4WtuVV5nladTv/rqd3zD2wGpLdijSXnvlYssRbSvR26fHonwz9ZD
LKmbp9gq/8SH7BUdDxPHJy/u+iIx+HuPdEB8AgPBAlNFSnoH9TklXqJf8IC1jnT9FDGjc3xSd6TT
FmadhiPHLzgjAN9pJwvNu89xE+PIs8m9lDONUe9mDInRPO+rCWMo3u7XRXNnOAZo7napqODnKNre
SJA/ELZVIwBdTEqwMLRMayQA7cSkutjGl5pBDRfeAZI+/e4GE4w3U8wHfXTCeRKx7dL0SdjDyW/C
mTDSgMJVfRO/bCuXG6RIKFg1bnWn5Xll8l7f+PHym3KtYTqokffe9iv/FP5hel0nYr44qm8/YhOI
EisM3zE9zpXnmSMnnWIZKDXxo3dECHlHJUu2qgINGOBdT6F/4/NSyWWnf4vrS/CTbboQGdxI1eE6
5gF+7aL/kLPoLNZMbTxWrA31NYgYy536ZIY4SjsBrAJsQSc76wQPHFQtO/z/vUo3mgti5MZwWprd
3IsrJa6gu+phS5PeFMd2XC43BVYHRL3xyBpvrtWRpVQdvLF0Y0f67j2/IF7YbqKFHbly/ZlfTpod
HV9LjjEBr4LPWlzz5l1oaFI2c8SAzSSjqSupeO2M3xQZJxW8UFtsAoThLOPc9jxAXV83AoSe9Qx3
TAt4QdxVIuGUiu8N7fArFLIFRu8xDlRY8sF64FqvQDkzbd99HCp4DmFKjyOLxolyTv6SBwnNaSgP
55P8W64Z3ZJG/f07vxy+6zPky5MG/HSYV4KPZVGKx5+FbI91RC7BjyqAGL8s674AmAmogunyMBEC
/hwwB64zcg2r+3MgHwYSs6Ql1HzArwtpbKLk2xMaQ5DbdQYJQUj62vIJF8loCHq0/ePgvz9SjSqi
n9i92T/A/YWHKN/LBh9xwGPiZqIXn2WOpUctlARw50Uuv98OJCqsAQ3JEv1c8Pac65StmEaZEQOd
DlyWFFdWznuqUWwfS7KZFlRiQ7xhbfVZ2ed3Xaao+Iwm0f40ziaT6NKNXUnQFSmcaR5I9Ca5glSG
YBsfm1Ts3hqjBY7XkFCm0nPhmj6xy+QCad5kKlW1keYgxlXU2JpUOe2e7p1yuQRMc19EG9eMkWOD
+AznNI5Yrgd8MqOsPtSlViapjk3VSRGFfRj1c3IAbYjb7Iw33Rk5BoMtL5jL3c+oN41YPMREEWT1
uIhcQ9GweWvSIq/w2vdtDyApqTWizZ29EYMcDs8m56EXbefjLlUpeYkKYv7TSefKhP3bOyuO2/fj
3lSEkg+8VhJCUHoQVG9VE5g48Mz8voTnj8CPmZDb4rNYmghqjiNDHnWFErCDlEAxRsOtJabDxSTf
bJGX4EcFV9gLMamuiWbBh+18bHXSivQdQcdCUhxP+k3JSrBNrHHr6OqTy1OirV9/fjK+3IWzuvwR
0BLIrEu9+DrZ2Q+AAdCaPI4LOv2UYS9Xw6TTi4AUcf45F15koYrt5uj7+rXQiGqmDkuhlgfmj7VJ
KmGnk6h/sweZafw=
`protect end_protected
